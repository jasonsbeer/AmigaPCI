-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 6 2024 13:45:26

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    TSn : in std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    LDSn : out std_logic;
    CASUn : in std_logic;
    RAS1n : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    DBRn : in std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RAMENn : out std_logic;
    RASn : out std_logic;
    TACKn : out std_logic;
    CLKEN : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10038\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9633\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9615\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9060\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9030\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8900\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8487\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8288\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8276\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8235\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7938\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7868\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7850\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7796\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7434\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7391\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7068\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6993\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6656\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6542\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6437\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4440\ : std_logic;
signal \N__4437\ : std_logic;
signal \N__4434\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4395\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4353\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4257\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4211\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4077\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4017\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3987\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3945\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3735\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3720\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK40_OUT_i_i\ : std_logic;
signal \CLK80_OUT_i_i\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.REG_TACK_7_0_cascade_\ : std_logic;
signal \U712_REG_SM.un1_STATE_COUNT_5_0_1\ : std_logic;
signal \U712_REG_SM.N_183_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_6\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.N_162_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_166_0\ : std_logic;
signal \C3_c\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_REG_SM.N_162_0\ : std_logic;
signal \U712_REG_SM.N_171_0_cascade_\ : std_logic;
signal \U712_REG_SM.RnW_m\ : std_logic;
signal \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_\ : std_logic;
signal \U712_REG_SM.N_165_0\ : std_logic;
signal \U712_REG_SM.N_167_0_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_167_0\ : std_logic;
signal \U712_REG_SM.N_176_0_cascade_\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_157_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_157_0_cascade_\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_176_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_5\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_192\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U712_REG_SM.N_171_0\ : std_logic;
signal \U712_REG_SM.UDS_OUT_2_0_0\ : std_logic;
signal \U712_REG_SM.LDS_OUTZ0\ : std_logic;
signal \U712_REG_SM_un1_LDSn_i\ : std_logic;
signal \U712_REG_SM.UDS_OUTZ0\ : std_logic;
signal \U712_REG_SM.DS_ENZ0\ : std_logic;
signal \U712_REG_SM_un1_UDSn_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_REG_SM.N_163_0\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_186\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_188\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_cascade_\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \U712_REG_SM.DS_EN_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_0\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \CLK40_OUT_i\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_CYCLE_TERM.N_45_0_0_en_0\ : std_logic;
signal \U712_REG_SM.LDS_OUT_2_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \N_614_i\ : std_logic;
signal \U712_CHIP_RAM.N_36\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \bfn_10_7_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.N_49_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_1\ : std_logic;
signal \U712_REG_SM_DBR_SYNC_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.N_57_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_58_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_40_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_99_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_85\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_65_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_58\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_0\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0_0_tz\ : std_logic;
signal \U712_BYTE_ENABLE.LW_TRANS_0\ : std_logic;
signal \U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_\ : std_logic;
signal \A_c_1\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U712_CHIP_RAM.N_34\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.N_74_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_50_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_75\ : std_logic;
signal \U712_CHIP_RAM.N_60\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_77\ : std_logic;
signal \U712_CHIP_RAM.N_40\ : std_logic;
signal \U712_CHIP_RAM.N_62_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_13_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_44_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_93\ : std_logic;
signal \U712_CHIP_RAM.N_13\ : std_logic;
signal \U712_CHIP_RAM.N_65\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_62\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_57\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CLLBEnZ0\ : std_logic;
signal \CLLBEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_38\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_6\ : std_logic;
signal \U712_CHIP_RAM.N_44\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.N_47\ : std_logic;
signal \U712_CHIP_RAM.N_47_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_89\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0\ : std_logic;
signal \U712_CHIP_RAM.N_100\ : std_logic;
signal \U712_CHIP_RAM.N_100_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_101\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_56\ : std_logic;
signal \U712_CHIP_RAM.N_42\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.N_42_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.N_98\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DRDDIR_0_i\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\ : std_logic;
signal \U712_CHIP_RAM.N_45\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\ : std_logic;
signal \A_c_18\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U712_CHIP_RAM.N_35\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_3\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_33\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_32\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CUMBEnZ0\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CUMBEn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CLMBEnZ0\ : std_logic;
signal \CLMBEn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.un2_CUUBEnZ0\ : std_logic;
signal \CUUBEn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \N_52_i\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.N_37\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.N_39\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \RASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA31_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_1\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \RAS1n_c\ : std_logic;
signal \U712_CHIP_RAM.RAS_SYNCZ0Z_0\ : std_logic;
signal \_gnd_net_\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \CLKEN_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \RAS0n_wire\ : std_logic;
signal \RAS1n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    CLKEN <= \CLKEN_wire\;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \RAS0n_wire\ <= RAS0n;
    \RAS1n_wire\ <= RAS1n;
    CMA <= \CMA_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    LDSn <= \LDSn_wire\;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_OUT_i\,
            REFERENCECLK => \N__3518\,
            RESETB => \N__8215\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_OUT\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10065\,
            DIN => \N__10064\,
            DOUT => \N__10063\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10065\,
            PADOUT => \N__10064\,
            PADIN => \N__10063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7598\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10056\,
            DIN => \N__10055\,
            DOUT => \N__10054\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10056\,
            PADOUT => \N__10055\,
            PADIN => \N__10054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10047\,
            DIN => \N__10046\,
            DOUT => \N__10045\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10047\,
            PADOUT => \N__10046\,
            PADIN => \N__10045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7979\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10038\,
            DIN => \N__10037\,
            DOUT => \N__10036\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10038\,
            PADOUT => \N__10037\,
            PADIN => \N__10036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10029\,
            DIN => \N__10028\,
            DOUT => \N__10027\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10029\,
            PADOUT => \N__10028\,
            PADIN => \N__10027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10020\,
            DIN => \N__10019\,
            DOUT => \N__10018\,
            PACKAGEPIN => \CLKEN_wire\
        );

    \CLKEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10020\,
            PADOUT => \N__10019\,
            PADIN => \N__10018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8219\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10011\,
            DIN => \N__10010\,
            DOUT => \N__10009\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__10011\,
            PADOUT => \N__10010\,
            PADIN => \N__10009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10002\,
            DIN => \N__10001\,
            DOUT => \N__10000\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10002\,
            PADOUT => \N__10001\,
            PADIN => \N__10000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9993\,
            DIN => \N__9992\,
            DOUT => \N__9991\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9993\,
            PADOUT => \N__9992\,
            PADIN => \N__9991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS1n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9984\,
            DIN => \N__9983\,
            DOUT => \N__9982\,
            PACKAGEPIN => \RAS1n_wire\
        );

    \RAS1n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9984\,
            PADOUT => \N__9983\,
            PADIN => \N__9982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS1n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9975\,
            DIN => \N__9974\,
            DOUT => \N__9973\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9975\,
            PADOUT => \N__9974\,
            PADIN => \N__9973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9966\,
            DIN => \N__9965\,
            DOUT => \N__9964\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9966\,
            PADOUT => \N__9965\,
            PADIN => \N__9964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7313\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9957\,
            DIN => \N__9956\,
            DOUT => \N__9955\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9957\,
            PADOUT => \N__9956\,
            PADIN => \N__9955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4942\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9948\,
            DIN => \N__9947\,
            DOUT => \N__9946\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9948\,
            PADOUT => \N__9947\,
            PADIN => \N__9946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9939\,
            DIN => \N__9938\,
            DOUT => \N__9937\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9939\,
            PADOUT => \N__9938\,
            PADIN => \N__9937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9930\,
            DIN => \N__9929\,
            DOUT => \N__9928\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9930\,
            PADOUT => \N__9929\,
            PADIN => \N__9928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9921\,
            DIN => \N__9920\,
            DOUT => \N__9919\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9921\,
            PADOUT => \N__9920\,
            PADIN => \N__9919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9912\,
            DIN => \N__9911\,
            DOUT => \N__9910\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9912\,
            PADOUT => \N__9911\,
            PADIN => \N__9910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9903\,
            DIN => \N__9902\,
            DOUT => \N__9901\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9903\,
            PADOUT => \N__9902\,
            PADIN => \N__9901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6899\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9894\,
            DIN => \N__9893\,
            DOUT => \N__9892\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9894\,
            PADOUT => \N__9893\,
            PADIN => \N__9892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9885\,
            DIN => \N__9884\,
            DOUT => \N__9883\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9885\,
            PADOUT => \N__9884\,
            PADIN => \N__9883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6542\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9876\,
            DIN => \N__9875\,
            DOUT => \N__9874\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9876\,
            PADOUT => \N__9875\,
            PADIN => \N__9874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9867\,
            DIN => \N__9866\,
            DOUT => \N__9865\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9867\,
            PADOUT => \N__9866\,
            PADIN => \N__9865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9858\,
            DIN => \N__9857\,
            DOUT => \N__9856\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9858\,
            PADOUT => \N__9857\,
            PADIN => \N__9856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9849\,
            DIN => \N__9848\,
            DOUT => \N__9847\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9849\,
            PADOUT => \N__9848\,
            PADIN => \N__9847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9840\,
            DIN => \N__9839\,
            DOUT => \N__9838\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9840\,
            PADOUT => \N__9839\,
            PADIN => \N__9838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9831\,
            DIN => \N__9830\,
            DOUT => \N__9829\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9831\,
            PADOUT => \N__9830\,
            PADIN => \N__9829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9822\,
            DIN => \N__9821\,
            DOUT => \N__9820\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9822\,
            PADOUT => \N__9821\,
            PADIN => \N__9820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9813\,
            DIN => \N__9812\,
            DOUT => \N__9811\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9813\,
            PADOUT => \N__9812\,
            PADIN => \N__9811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9804\,
            DIN => \N__9803\,
            DOUT => \N__9802\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9804\,
            PADOUT => \N__9803\,
            PADIN => \N__9802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9795\,
            DIN => \N__9794\,
            DOUT => \N__9793\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9795\,
            PADOUT => \N__9794\,
            PADIN => \N__9793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9786\,
            DIN => \N__9785\,
            DOUT => \N__9784\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9786\,
            PADOUT => \N__9785\,
            PADIN => \N__9784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5501\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9777\,
            DIN => \N__9776\,
            DOUT => \N__9775\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9777\,
            PADOUT => \N__9776\,
            PADIN => \N__9775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9768\,
            DIN => \N__9767\,
            DOUT => \N__9766\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9768\,
            PADOUT => \N__9767\,
            PADIN => \N__9766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9759\,
            DIN => \N__9758\,
            DOUT => \N__9757\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9759\,
            PADOUT => \N__9758\,
            PADIN => \N__9757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9750\,
            DIN => \N__9749\,
            DOUT => \N__9748\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9750\,
            PADOUT => \N__9749\,
            PADIN => \N__9748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9741\,
            DIN => \N__9740\,
            DOUT => \N__9739\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9741\,
            PADOUT => \N__9740\,
            PADIN => \N__9739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9732\,
            DIN => \N__9731\,
            DOUT => \N__9730\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9732\,
            PADOUT => \N__9731\,
            PADIN => \N__9730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9723\,
            DIN => \N__9722\,
            DOUT => \N__9721\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9723\,
            PADOUT => \N__9722\,
            PADIN => \N__9721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9714\,
            DIN => \N__9713\,
            DOUT => \N__9712\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9714\,
            PADOUT => \N__9713\,
            PADIN => \N__9712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7679\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9705\,
            DIN => \N__9704\,
            DOUT => \N__9703\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9705\,
            PADOUT => \N__9704\,
            PADIN => \N__9703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9696\,
            DIN => \N__9695\,
            DOUT => \N__9694\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9696\,
            PADOUT => \N__9695\,
            PADIN => \N__9694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9687\,
            DIN => \N__9686\,
            DOUT => \N__9685\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9687\,
            PADOUT => \N__9686\,
            PADIN => \N__9685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3584\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9678\,
            DIN => \N__9677\,
            DOUT => \N__9676\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9678\,
            PADOUT => \N__9677\,
            PADIN => \N__9676\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9669\,
            DIN => \N__9668\,
            DOUT => \N__9667\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9669\,
            PADOUT => \N__9668\,
            PADIN => \N__9667\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3566\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9660\,
            DIN => \N__9659\,
            DOUT => \N__9658\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9660\,
            PADOUT => \N__9659\,
            PADIN => \N__9658\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6881\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9651\,
            DIN => \N__9650\,
            DOUT => \N__9649\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9651\,
            PADOUT => \N__9650\,
            PADIN => \N__9649\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9642\,
            DIN => \N__9641\,
            DOUT => \N__9640\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9642\,
            PADOUT => \N__9641\,
            PADIN => \N__9640\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9633\,
            DIN => \N__9632\,
            DOUT => \N__9631\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9633\,
            PADOUT => \N__9632\,
            PADIN => \N__9631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9624\,
            DIN => \N__9623\,
            DOUT => \N__9622\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9624\,
            PADOUT => \N__9623\,
            PADIN => \N__9622\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9615\,
            DIN => \N__9614\,
            DOUT => \N__9613\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9615\,
            PADOUT => \N__9614\,
            PADIN => \N__9613\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9606\,
            DIN => \N__9605\,
            DOUT => \N__9604\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9606\,
            PADOUT => \N__9605\,
            PADIN => \N__9604\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4571\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9597\,
            DIN => \N__9596\,
            DOUT => \N__9595\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9597\,
            PADOUT => \N__9596\,
            PADIN => \N__9595\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7406\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9588\,
            DIN => \N__9587\,
            DOUT => \N__9586\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9588\,
            PADOUT => \N__9587\,
            PADIN => \N__9586\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9579\,
            DIN => \N__9578\,
            DOUT => \N__9577\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9579\,
            PADOUT => \N__9578\,
            PADIN => \N__9577\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7271\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9570\,
            DIN => \N__9569\,
            DOUT => \N__9568\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9570\,
            PADOUT => \N__9569\,
            PADIN => \N__9568\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3562\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9561\,
            DIN => \N__9560\,
            DOUT => \N__9559\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9561\,
            PADOUT => \N__9560\,
            PADIN => \N__9559\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9552\,
            DIN => \N__9551\,
            DOUT => \N__9550\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9552\,
            PADOUT => \N__9551\,
            PADIN => \N__9550\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9543\,
            DIN => \N__9542\,
            DOUT => \N__9541\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9543\,
            PADOUT => \N__9542\,
            PADIN => \N__9541\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9534\,
            DIN => \N__9533\,
            DOUT => \N__9532\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9534\,
            PADOUT => \N__9533\,
            PADIN => \N__9532\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8897\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9525\,
            DIN => \N__9524\,
            DOUT => \N__9523\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9525\,
            PADOUT => \N__9524\,
            PADIN => \N__9523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6695\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9516\,
            DIN => \N__9515\,
            DOUT => \N__9514\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9516\,
            PADOUT => \N__9515\,
            PADIN => \N__9514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9507\,
            DIN => \N__9506\,
            DOUT => \N__9505\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9507\,
            PADOUT => \N__9506\,
            PADIN => \N__9505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9498\,
            DIN => \N__9497\,
            DOUT => \N__9496\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9498\,
            PADOUT => \N__9497\,
            PADIN => \N__9496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9489\,
            DIN => \N__9488\,
            DOUT => \N__9487\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9489\,
            PADOUT => \N__9488\,
            PADIN => \N__9487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9480\,
            DIN => \N__9479\,
            DOUT => \N__9478\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9480\,
            PADOUT => \N__9479\,
            PADIN => \N__9478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9471\,
            DIN => \N__9470\,
            DOUT => \N__9469\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9471\,
            PADOUT => \N__9470\,
            PADIN => \N__9469\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6464\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9462\,
            DIN => \N__9461\,
            DOUT => \N__9460\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9462\,
            PADOUT => \N__9461\,
            PADIN => \N__9460\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9453\,
            DIN => \N__9452\,
            DOUT => \N__9451\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9453\,
            PADOUT => \N__9452\,
            PADIN => \N__9451\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7532\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9444\,
            DIN => \N__9443\,
            DOUT => \N__9442\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__9444\,
            PADOUT => \N__9443\,
            PADIN => \N__9442\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4598\,
            DIN0 => OPEN,
            DOUT0 => \N__3842\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9435\,
            DIN => \N__9434\,
            DOUT => \N__9433\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9435\,
            PADOUT => \N__9434\,
            PADIN => \N__9433\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9426\,
            DIN => \N__9425\,
            DOUT => \N__9424\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9426\,
            PADOUT => \N__9425\,
            PADIN => \N__9424\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9417\,
            DIN => \N__9416\,
            DOUT => \N__9415\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9417\,
            PADOUT => \N__9416\,
            PADIN => \N__9415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9408\,
            DIN => \N__9407\,
            DOUT => \N__9406\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9408\,
            PADOUT => \N__9407\,
            PADIN => \N__9406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8675\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9399\,
            DIN => \N__9398\,
            DOUT => \N__9397\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9399\,
            PADOUT => \N__9398\,
            PADIN => \N__9397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9390\,
            DIN => \N__9389\,
            DOUT => \N__9388\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9390\,
            PADOUT => \N__9389\,
            PADIN => \N__9388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9381\,
            DIN => \N__9380\,
            DOUT => \N__9379\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9381\,
            PADOUT => \N__9380\,
            PADIN => \N__9379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9372\,
            DIN => \N__9371\,
            DOUT => \N__9370\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9372\,
            PADOUT => \N__9371\,
            PADIN => \N__9370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9363\,
            DIN => \N__9362\,
            DOUT => \N__9361\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9363\,
            PADOUT => \N__9362\,
            PADIN => \N__9361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9354\,
            DIN => \N__9353\,
            DOUT => \N__9352\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9354\,
            PADOUT => \N__9353\,
            PADIN => \N__9352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4244\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2241\ : CascadeMux
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9329\,
            I => \N__9325\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__2237\ : Span4Mux_h
    port map (
            O => \N__9325\,
            I => \N__9317\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9322\,
            I => \N__9317\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__9317\,
            I => \N__9314\
        );

    \I__2234\ : Sp12to4
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__2233\ : Odrv12
    port map (
            O => \N__9311\,
            I => \RAS0n_c\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9305\,
            I => \N__9302\
        );

    \I__2230\ : Odrv12
    port map (
            O => \N__9302\,
            I => \RAS1n_c\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9299\,
            I => \N__9295\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9292\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9295\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9292\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9287\,
            I => \N__9284\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9284\,
            I => \N__9242\
        );

    \I__2223\ : ClkMux
    port map (
            O => \N__9283\,
            I => \N__9125\
        );

    \I__2222\ : ClkMux
    port map (
            O => \N__9282\,
            I => \N__9125\
        );

    \I__2221\ : ClkMux
    port map (
            O => \N__9281\,
            I => \N__9125\
        );

    \I__2220\ : ClkMux
    port map (
            O => \N__9280\,
            I => \N__9125\
        );

    \I__2219\ : ClkMux
    port map (
            O => \N__9279\,
            I => \N__9125\
        );

    \I__2218\ : ClkMux
    port map (
            O => \N__9278\,
            I => \N__9125\
        );

    \I__2217\ : ClkMux
    port map (
            O => \N__9277\,
            I => \N__9125\
        );

    \I__2216\ : ClkMux
    port map (
            O => \N__9276\,
            I => \N__9125\
        );

    \I__2215\ : ClkMux
    port map (
            O => \N__9275\,
            I => \N__9125\
        );

    \I__2214\ : ClkMux
    port map (
            O => \N__9274\,
            I => \N__9125\
        );

    \I__2213\ : ClkMux
    port map (
            O => \N__9273\,
            I => \N__9125\
        );

    \I__2212\ : ClkMux
    port map (
            O => \N__9272\,
            I => \N__9125\
        );

    \I__2211\ : ClkMux
    port map (
            O => \N__9271\,
            I => \N__9125\
        );

    \I__2210\ : ClkMux
    port map (
            O => \N__9270\,
            I => \N__9125\
        );

    \I__2209\ : ClkMux
    port map (
            O => \N__9269\,
            I => \N__9125\
        );

    \I__2208\ : ClkMux
    port map (
            O => \N__9268\,
            I => \N__9125\
        );

    \I__2207\ : ClkMux
    port map (
            O => \N__9267\,
            I => \N__9125\
        );

    \I__2206\ : ClkMux
    port map (
            O => \N__9266\,
            I => \N__9125\
        );

    \I__2205\ : ClkMux
    port map (
            O => \N__9265\,
            I => \N__9125\
        );

    \I__2204\ : ClkMux
    port map (
            O => \N__9264\,
            I => \N__9125\
        );

    \I__2203\ : ClkMux
    port map (
            O => \N__9263\,
            I => \N__9125\
        );

    \I__2202\ : ClkMux
    port map (
            O => \N__9262\,
            I => \N__9125\
        );

    \I__2201\ : ClkMux
    port map (
            O => \N__9261\,
            I => \N__9125\
        );

    \I__2200\ : ClkMux
    port map (
            O => \N__9260\,
            I => \N__9125\
        );

    \I__2199\ : ClkMux
    port map (
            O => \N__9259\,
            I => \N__9125\
        );

    \I__2198\ : ClkMux
    port map (
            O => \N__9258\,
            I => \N__9125\
        );

    \I__2197\ : ClkMux
    port map (
            O => \N__9257\,
            I => \N__9125\
        );

    \I__2196\ : ClkMux
    port map (
            O => \N__9256\,
            I => \N__9125\
        );

    \I__2195\ : ClkMux
    port map (
            O => \N__9255\,
            I => \N__9125\
        );

    \I__2194\ : ClkMux
    port map (
            O => \N__9254\,
            I => \N__9125\
        );

    \I__2193\ : ClkMux
    port map (
            O => \N__9253\,
            I => \N__9125\
        );

    \I__2192\ : ClkMux
    port map (
            O => \N__9252\,
            I => \N__9125\
        );

    \I__2191\ : ClkMux
    port map (
            O => \N__9251\,
            I => \N__9125\
        );

    \I__2190\ : ClkMux
    port map (
            O => \N__9250\,
            I => \N__9125\
        );

    \I__2189\ : ClkMux
    port map (
            O => \N__9249\,
            I => \N__9125\
        );

    \I__2188\ : ClkMux
    port map (
            O => \N__9248\,
            I => \N__9125\
        );

    \I__2187\ : ClkMux
    port map (
            O => \N__9247\,
            I => \N__9125\
        );

    \I__2186\ : ClkMux
    port map (
            O => \N__9246\,
            I => \N__9125\
        );

    \I__2185\ : ClkMux
    port map (
            O => \N__9245\,
            I => \N__9125\
        );

    \I__2184\ : Glb2LocalMux
    port map (
            O => \N__9242\,
            I => \N__9125\
        );

    \I__2183\ : ClkMux
    port map (
            O => \N__9241\,
            I => \N__9125\
        );

    \I__2182\ : ClkMux
    port map (
            O => \N__9240\,
            I => \N__9125\
        );

    \I__2181\ : ClkMux
    port map (
            O => \N__9239\,
            I => \N__9125\
        );

    \I__2180\ : ClkMux
    port map (
            O => \N__9238\,
            I => \N__9125\
        );

    \I__2179\ : ClkMux
    port map (
            O => \N__9237\,
            I => \N__9125\
        );

    \I__2178\ : ClkMux
    port map (
            O => \N__9236\,
            I => \N__9125\
        );

    \I__2177\ : ClkMux
    port map (
            O => \N__9235\,
            I => \N__9125\
        );

    \I__2176\ : ClkMux
    port map (
            O => \N__9234\,
            I => \N__9125\
        );

    \I__2175\ : ClkMux
    port map (
            O => \N__9233\,
            I => \N__9125\
        );

    \I__2174\ : ClkMux
    port map (
            O => \N__9232\,
            I => \N__9125\
        );

    \I__2173\ : ClkMux
    port map (
            O => \N__9231\,
            I => \N__9125\
        );

    \I__2172\ : ClkMux
    port map (
            O => \N__9230\,
            I => \N__9125\
        );

    \I__2171\ : GlobalMux
    port map (
            O => \N__9125\,
            I => \CLK80_OUT\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9113\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9107\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9104\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9101\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9098\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9095\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9092\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9085\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9085\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9085\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9082\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9073\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9048\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__9101\,
            I => \N__9045\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9098\,
            I => \N__9038\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9095\,
            I => \N__9030\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9092\,
            I => \N__9027\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9085\,
            I => \N__9019\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9015\
        );

    \I__2151\ : SRMux
    port map (
            O => \N__9081\,
            I => \N__8903\
        );

    \I__2150\ : SRMux
    port map (
            O => \N__9080\,
            I => \N__8903\
        );

    \I__2149\ : SRMux
    port map (
            O => \N__9079\,
            I => \N__8903\
        );

    \I__2148\ : SRMux
    port map (
            O => \N__9078\,
            I => \N__8903\
        );

    \I__2147\ : SRMux
    port map (
            O => \N__9077\,
            I => \N__8903\
        );

    \I__2146\ : SRMux
    port map (
            O => \N__9076\,
            I => \N__8903\
        );

    \I__2145\ : Glb2LocalMux
    port map (
            O => \N__9073\,
            I => \N__8903\
        );

    \I__2144\ : SRMux
    port map (
            O => \N__9072\,
            I => \N__8903\
        );

    \I__2143\ : SRMux
    port map (
            O => \N__9071\,
            I => \N__8903\
        );

    \I__2142\ : SRMux
    port map (
            O => \N__9070\,
            I => \N__8903\
        );

    \I__2141\ : SRMux
    port map (
            O => \N__9069\,
            I => \N__8903\
        );

    \I__2140\ : SRMux
    port map (
            O => \N__9068\,
            I => \N__8903\
        );

    \I__2139\ : SRMux
    port map (
            O => \N__9067\,
            I => \N__8903\
        );

    \I__2138\ : SRMux
    port map (
            O => \N__9066\,
            I => \N__8903\
        );

    \I__2137\ : SRMux
    port map (
            O => \N__9065\,
            I => \N__8903\
        );

    \I__2136\ : SRMux
    port map (
            O => \N__9064\,
            I => \N__8903\
        );

    \I__2135\ : SRMux
    port map (
            O => \N__9063\,
            I => \N__8903\
        );

    \I__2134\ : SRMux
    port map (
            O => \N__9062\,
            I => \N__8903\
        );

    \I__2133\ : SRMux
    port map (
            O => \N__9061\,
            I => \N__8903\
        );

    \I__2132\ : SRMux
    port map (
            O => \N__9060\,
            I => \N__8903\
        );

    \I__2131\ : SRMux
    port map (
            O => \N__9059\,
            I => \N__8903\
        );

    \I__2130\ : SRMux
    port map (
            O => \N__9058\,
            I => \N__8903\
        );

    \I__2129\ : SRMux
    port map (
            O => \N__9057\,
            I => \N__8903\
        );

    \I__2128\ : SRMux
    port map (
            O => \N__9056\,
            I => \N__8903\
        );

    \I__2127\ : SRMux
    port map (
            O => \N__9055\,
            I => \N__8903\
        );

    \I__2126\ : SRMux
    port map (
            O => \N__9054\,
            I => \N__8903\
        );

    \I__2125\ : SRMux
    port map (
            O => \N__9053\,
            I => \N__8903\
        );

    \I__2124\ : SRMux
    port map (
            O => \N__9052\,
            I => \N__8903\
        );

    \I__2123\ : SRMux
    port map (
            O => \N__9051\,
            I => \N__8903\
        );

    \I__2122\ : Glb2LocalMux
    port map (
            O => \N__9048\,
            I => \N__8903\
        );

    \I__2121\ : Glb2LocalMux
    port map (
            O => \N__9045\,
            I => \N__8903\
        );

    \I__2120\ : SRMux
    port map (
            O => \N__9044\,
            I => \N__8903\
        );

    \I__2119\ : SRMux
    port map (
            O => \N__9043\,
            I => \N__8903\
        );

    \I__2118\ : SRMux
    port map (
            O => \N__9042\,
            I => \N__8903\
        );

    \I__2117\ : SRMux
    port map (
            O => \N__9041\,
            I => \N__8903\
        );

    \I__2116\ : Glb2LocalMux
    port map (
            O => \N__9038\,
            I => \N__8903\
        );

    \I__2115\ : SRMux
    port map (
            O => \N__9037\,
            I => \N__8903\
        );

    \I__2114\ : SRMux
    port map (
            O => \N__9036\,
            I => \N__8903\
        );

    \I__2113\ : SRMux
    port map (
            O => \N__9035\,
            I => \N__8903\
        );

    \I__2112\ : SRMux
    port map (
            O => \N__9034\,
            I => \N__8903\
        );

    \I__2111\ : SRMux
    port map (
            O => \N__9033\,
            I => \N__8903\
        );

    \I__2110\ : Glb2LocalMux
    port map (
            O => \N__9030\,
            I => \N__8903\
        );

    \I__2109\ : Glb2LocalMux
    port map (
            O => \N__9027\,
            I => \N__8903\
        );

    \I__2108\ : SRMux
    port map (
            O => \N__9026\,
            I => \N__8903\
        );

    \I__2107\ : SRMux
    port map (
            O => \N__9025\,
            I => \N__8903\
        );

    \I__2106\ : SRMux
    port map (
            O => \N__9024\,
            I => \N__8903\
        );

    \I__2105\ : SRMux
    port map (
            O => \N__9023\,
            I => \N__8903\
        );

    \I__2104\ : SRMux
    port map (
            O => \N__9022\,
            I => \N__8903\
        );

    \I__2103\ : Glb2LocalMux
    port map (
            O => \N__9019\,
            I => \N__8903\
        );

    \I__2102\ : SRMux
    port map (
            O => \N__9018\,
            I => \N__8903\
        );

    \I__2101\ : Glb2LocalMux
    port map (
            O => \N__9015\,
            I => \N__8903\
        );

    \I__2100\ : SRMux
    port map (
            O => \N__9014\,
            I => \N__8903\
        );

    \I__2099\ : SRMux
    port map (
            O => \N__9013\,
            I => \N__8903\
        );

    \I__2098\ : SRMux
    port map (
            O => \N__9012\,
            I => \N__8903\
        );

    \I__2097\ : GlobalMux
    port map (
            O => \N__8903\,
            I => \N__8900\
        );

    \I__2096\ : gio2CtrlBuf
    port map (
            O => \N__8900\,
            I => \RESETn_c_i_g\
        );

    \I__2095\ : IoInMux
    port map (
            O => \N__8897\,
            I => \N__8894\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__8894\,
            I => \N__8891\
        );

    \I__2093\ : Span4Mux_s2_h
    port map (
            O => \N__8891\,
            I => \N__8888\
        );

    \I__2092\ : Sp12to4
    port map (
            O => \N__8888\,
            I => \N__8885\
        );

    \I__2091\ : Span12Mux_s8_v
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__2090\ : Odrv12
    port map (
            O => \N__8882\,
            I => \WEn_c\
        );

    \I__2089\ : InMux
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__8876\,
            I => \N__8873\
        );

    \I__2087\ : Span12Mux_v
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__2086\ : Span12Mux_h
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__2085\ : Odrv12
    port map (
            O => \N__8867\,
            I => \A_c_17\
        );

    \I__2084\ : InMux
    port map (
            O => \N__8864\,
            I => \N__8858\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__8863\,
            I => \N__8853\
        );

    \I__2082\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8845\
        );

    \I__2081\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8835\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__8858\,
            I => \N__8832\
        );

    \I__2079\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8827\
        );

    \I__2078\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8827\
        );

    \I__2077\ : InMux
    port map (
            O => \N__8853\,
            I => \N__8819\
        );

    \I__2076\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8819\
        );

    \I__2075\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8819\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8816\
        );

    \I__2073\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8813\
        );

    \I__2072\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8810\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__8845\,
            I => \N__8807\
        );

    \I__2070\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8802\
        );

    \I__2069\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8802\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8797\
        );

    \I__2067\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8797\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8791\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8788\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8784\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8835\,
            I => \N__8777\
        );

    \I__2062\ : Span4Mux_v
    port map (
            O => \N__8832\,
            I => \N__8777\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__8827\,
            I => \N__8777\
        );

    \I__2060\ : InMux
    port map (
            O => \N__8826\,
            I => \N__8774\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8769\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__8816\,
            I => \N__8769\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8813\,
            I => \N__8761\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__8810\,
            I => \N__8758\
        );

    \I__2055\ : Span4Mux_v
    port map (
            O => \N__8807\,
            I => \N__8755\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__8802\,
            I => \N__8750\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8750\
        );

    \I__2052\ : InMux
    port map (
            O => \N__8796\,
            I => \N__8745\
        );

    \I__2051\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8745\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8742\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__8791\,
            I => \N__8737\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__8788\,
            I => \N__8737\
        );

    \I__2047\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8734\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__8784\,
            I => \N__8727\
        );

    \I__2045\ : Span4Mux_v
    port map (
            O => \N__8777\,
            I => \N__8727\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__8774\,
            I => \N__8727\
        );

    \I__2043\ : Span4Mux_v
    port map (
            O => \N__8769\,
            I => \N__8724\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8721\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8718\
        );

    \I__2040\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8711\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8711\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8711\
        );

    \I__2037\ : Span4Mux_v
    port map (
            O => \N__8761\,
            I => \N__8704\
        );

    \I__2036\ : Span4Mux_h
    port map (
            O => \N__8758\,
            I => \N__8704\
        );

    \I__2035\ : Span4Mux_v
    port map (
            O => \N__8755\,
            I => \N__8704\
        );

    \I__2034\ : Span4Mux_v
    port map (
            O => \N__8750\,
            I => \N__8699\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8699\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8742\,
            I => \N__8690\
        );

    \I__2031\ : Span4Mux_h
    port map (
            O => \N__8737\,
            I => \N__8690\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__8734\,
            I => \N__8690\
        );

    \I__2029\ : Span4Mux_h
    port map (
            O => \N__8727\,
            I => \N__8690\
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__8724\,
            I => \CPU_CYCLEm\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8721\,
            I => \CPU_CYCLEm\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8718\,
            I => \CPU_CYCLEm\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8711\,
            I => \CPU_CYCLEm\
        );

    \I__2024\ : Odrv4
    port map (
            O => \N__8704\,
            I => \CPU_CYCLEm\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__8699\,
            I => \CPU_CYCLEm\
        );

    \I__2022\ : Odrv4
    port map (
            O => \N__8690\,
            I => \CPU_CYCLEm\
        );

    \I__2021\ : IoInMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__2019\ : IoSpan4Mux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__2018\ : Span4Mux_s3_h
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__2015\ : Odrv4
    port map (
            O => \N__8657\,
            I => \CMA_c_8\
        );

    \I__2014\ : CEMux
    port map (
            O => \N__8654\,
            I => \N__8650\
        );

    \I__2013\ : CEMux
    port map (
            O => \N__8653\,
            I => \N__8647\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__8650\,
            I => \N__8640\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8647\,
            I => \N__8640\
        );

    \I__2010\ : CEMux
    port map (
            O => \N__8646\,
            I => \N__8637\
        );

    \I__2009\ : CEMux
    port map (
            O => \N__8645\,
            I => \N__8634\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__8640\,
            I => \N__8628\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8637\,
            I => \N__8628\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8634\,
            I => \N__8625\
        );

    \I__2005\ : CEMux
    port map (
            O => \N__8633\,
            I => \N__8622\
        );

    \I__2004\ : Span4Mux_h
    port map (
            O => \N__8628\,
            I => \N__8618\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__8625\,
            I => \N__8613\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8610\
        );

    \I__2001\ : CEMux
    port map (
            O => \N__8621\,
            I => \N__8607\
        );

    \I__2000\ : Span4Mux_h
    port map (
            O => \N__8618\,
            I => \N__8604\
        );

    \I__1999\ : CEMux
    port map (
            O => \N__8617\,
            I => \N__8601\
        );

    \I__1998\ : CEMux
    port map (
            O => \N__8616\,
            I => \N__8598\
        );

    \I__1997\ : Odrv4
    port map (
            O => \N__8613\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__8610\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8607\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__8604\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8601\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__8598\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i_0\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8578\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8569\
        );

    \I__1989\ : InMux
    port map (
            O => \N__8583\,
            I => \N__8569\
        );

    \I__1988\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8564\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8564\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8578\,
            I => \N__8561\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8558\
        );

    \I__1984\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8553\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8549\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8546\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8543\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8564\,
            I => \N__8538\
        );

    \I__1979\ : Span4Mux_h
    port map (
            O => \N__8561\,
            I => \N__8538\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8535\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__8557\,
            I => \N__8532\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8529\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8526\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8523\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__8549\,
            I => \N__8518\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8546\,
            I => \N__8518\
        );

    \I__1971\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8511\
        );

    \I__1970\ : Span4Mux_v
    port map (
            O => \N__8538\,
            I => \N__8511\
        );

    \I__1969\ : Span4Mux_h
    port map (
            O => \N__8535\,
            I => \N__8511\
        );

    \I__1968\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8506\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8503\
        );

    \I__1966\ : Span4Mux_v
    port map (
            O => \N__8526\,
            I => \N__8500\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8523\,
            I => \N__8495\
        );

    \I__1964\ : Span4Mux_h
    port map (
            O => \N__8518\,
            I => \N__8495\
        );

    \I__1963\ : Span4Mux_h
    port map (
            O => \N__8511\,
            I => \N__8492\
        );

    \I__1962\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8487\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8487\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8506\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__8503\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__8500\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1957\ : Odrv4
    port map (
            O => \N__8495\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__8492\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8487\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__8474\,
            I => \N__8467\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__8473\,
            I => \N__8464\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__8472\,
            I => \N__8458\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__8471\,
            I => \N__8455\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8470\,
            I => \N__8451\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8467\,
            I => \N__8446\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8446\
        );

    \I__1947\ : InMux
    port map (
            O => \N__8463\,
            I => \N__8443\
        );

    \I__1946\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8437\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8437\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8458\,
            I => \N__8434\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8430\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8427\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__8451\,
            I => \N__8424\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8446\,
            I => \N__8421\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__8443\,
            I => \N__8418\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8442\,
            I => \N__8413\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8410\
        );

    \I__1936\ : LocalMux
    port map (
            O => \N__8434\,
            I => \N__8407\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8404\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__8430\,
            I => \N__8401\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8398\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__8424\,
            I => \N__8395\
        );

    \I__1931\ : Span4Mux_v
    port map (
            O => \N__8421\,
            I => \N__8390\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__8418\,
            I => \N__8390\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \N__8386\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8416\,
            I => \N__8383\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8380\
        );

    \I__1926\ : Span4Mux_h
    port map (
            O => \N__8410\,
            I => \N__8375\
        );

    \I__1925\ : Span4Mux_h
    port map (
            O => \N__8407\,
            I => \N__8375\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8370\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__8401\,
            I => \N__8370\
        );

    \I__1922\ : Span4Mux_v
    port map (
            O => \N__8398\,
            I => \N__8365\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__8395\,
            I => \N__8365\
        );

    \I__1920\ : Span4Mux_h
    port map (
            O => \N__8390\,
            I => \N__8362\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8357\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8357\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8383\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1916\ : Odrv12
    port map (
            O => \N__8380\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1915\ : Odrv4
    port map (
            O => \N__8375\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1914\ : Odrv4
    port map (
            O => \N__8370\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__8365\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1912\ : Odrv4
    port map (
            O => \N__8362\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8357\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8338\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8338\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8335\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1906\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8327\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8327\,
            I => \N__8324\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__8324\,
            I => \N__8320\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__1902\ : Sp12to4
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__8317\,
            I => \N__8311\
        );

    \I__1900\ : Span12Mux_h
    port map (
            O => \N__8314\,
            I => \N__8308\
        );

    \I__1899\ : Span12Mux_v
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__1898\ : Span12Mux_v
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1897\ : Span12Mux_h
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1896\ : Odrv12
    port map (
            O => \N__8302\,
            I => \DRA_c_4\
        );

    \I__1895\ : Odrv12
    port map (
            O => \N__8299\,
            I => \DRA_c_4\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8294\,
            I => \N__8291\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__8291\,
            I => \N__8288\
        );

    \I__1892\ : Odrv4
    port map (
            O => \N__8288\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1891\ : CEMux
    port map (
            O => \N__8285\,
            I => \N__8282\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8282\,
            I => \N__8276\
        );

    \I__1889\ : CEMux
    port map (
            O => \N__8281\,
            I => \N__8273\
        );

    \I__1888\ : CEMux
    port map (
            O => \N__8280\,
            I => \N__8270\
        );

    \I__1887\ : CEMux
    port map (
            O => \N__8279\,
            I => \N__8267\
        );

    \I__1886\ : Span4Mux_h
    port map (
            O => \N__8276\,
            I => \N__8263\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8273\,
            I => \N__8258\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__8270\,
            I => \N__8258\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__8267\,
            I => \N__8255\
        );

    \I__1882\ : CEMux
    port map (
            O => \N__8266\,
            I => \N__8252\
        );

    \I__1881\ : Span4Mux_h
    port map (
            O => \N__8263\,
            I => \N__8247\
        );

    \I__1880\ : Span4Mux_h
    port map (
            O => \N__8258\,
            I => \N__8244\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__8255\,
            I => \N__8241\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8252\,
            I => \N__8238\
        );

    \I__1877\ : CEMux
    port map (
            O => \N__8251\,
            I => \N__8235\
        );

    \I__1876\ : CEMux
    port map (
            O => \N__8250\,
            I => \N__8232\
        );

    \I__1875\ : Odrv4
    port map (
            O => \N__8247\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__8244\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__8241\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1872\ : Odrv12
    port map (
            O => \N__8238\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8235\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8232\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\
        );

    \I__1869\ : IoInMux
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8212\
        );

    \I__1867\ : IoInMux
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__1866\ : IoSpan4Mux
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1864\ : IoSpan4Mux
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__1863\ : Span4Mux_s2_v
    port map (
            O => \N__8203\,
            I => \N__8197\
        );

    \I__1862\ : Span4Mux_s3_h
    port map (
            O => \N__8200\,
            I => \N__8194\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__8197\,
            I => \N__8191\
        );

    \I__1860\ : Span4Mux_h
    port map (
            O => \N__8194\,
            I => \N__8188\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__8191\,
            I => \N__8185\
        );

    \I__1858\ : Odrv4
    port map (
            O => \N__8188\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__8185\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8173\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8176\,
            I => \N__8170\
        );

    \I__1853\ : Span4Mux_v
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8170\,
            I => \N__8164\
        );

    \I__1851\ : Sp12to4
    port map (
            O => \N__8167\,
            I => \N__8161\
        );

    \I__1850\ : Span4Mux_v
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1849\ : Span12Mux_h
    port map (
            O => \N__8161\,
            I => \N__8155\
        );

    \I__1848\ : Sp12to4
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__1847\ : Odrv12
    port map (
            O => \N__8155\,
            I => \DRA_c_8\
        );

    \I__1846\ : Odrv12
    port map (
            O => \N__8152\,
            I => \DRA_c_8\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8138\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__8138\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8135\,
            I => \N__8130\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__8134\,
            I => \N__8126\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__8133\,
            I => \N__8120\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8130\,
            I => \N__8111\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8108\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8105\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__8125\,
            I => \N__8102\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__8124\,
            I => \N__8099\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8096\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8093\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8090\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8118\,
            I => \N__8087\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8117\,
            I => \N__8084\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__8116\,
            I => \N__8081\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__8115\,
            I => \N__8078\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__8114\,
            I => \N__8075\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8111\,
            I => \N__8072\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8108\,
            I => \N__8067\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8105\,
            I => \N__8067\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8102\,
            I => \N__8062\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8062\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8096\,
            I => \N__8057\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8054\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8090\,
            I => \N__8051\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8048\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8084\,
            I => \N__8045\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8042\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8078\,
            I => \N__8039\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8075\,
            I => \N__8036\
        );

    \I__1812\ : Span4Mux_h
    port map (
            O => \N__8072\,
            I => \N__8029\
        );

    \I__1811\ : Span4Mux_v
    port map (
            O => \N__8067\,
            I => \N__8029\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8029\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__8061\,
            I => \N__8026\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8022\
        );

    \I__1807\ : Span4Mux_v
    port map (
            O => \N__8057\,
            I => \N__8017\
        );

    \I__1806\ : Span4Mux_v
    port map (
            O => \N__8054\,
            I => \N__8017\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__8051\,
            I => \N__8012\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__8012\
        );

    \I__1803\ : Span12Mux_v
    port map (
            O => \N__8045\,
            I => \N__8005\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8042\,
            I => \N__8005\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8039\,
            I => \N__8005\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8036\,
            I => \N__8002\
        );

    \I__1799\ : Span4Mux_h
    port map (
            O => \N__8029\,
            I => \N__7999\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8026\,
            I => \N__7994\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8025\,
            I => \N__7994\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8022\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1795\ : Odrv4
    port map (
            O => \N__8017\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__8012\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1793\ : Odrv12
    port map (
            O => \N__8005\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__8002\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__7999\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__7994\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1789\ : IoInMux
    port map (
            O => \N__7979\,
            I => \N__7976\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7973\
        );

    \I__1787\ : IoSpan4Mux
    port map (
            O => \N__7973\,
            I => \N__7970\
        );

    \I__1786\ : Sp12to4
    port map (
            O => \N__7970\,
            I => \N__7967\
        );

    \I__1785\ : Span12Mux_s9_v
    port map (
            O => \N__7967\,
            I => \N__7964\
        );

    \I__1784\ : Odrv12
    port map (
            O => \N__7964\,
            I => \CASn_c\
        );

    \I__1783\ : CEMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7953\
        );

    \I__1781\ : CEMux
    port map (
            O => \N__7957\,
            I => \N__7950\
        );

    \I__1780\ : CEMux
    port map (
            O => \N__7956\,
            I => \N__7947\
        );

    \I__1779\ : Span4Mux_v
    port map (
            O => \N__7953\,
            I => \N__7942\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__7950\,
            I => \N__7942\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7947\,
            I => \N__7938\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__7942\,
            I => \N__7935\
        );

    \I__1775\ : CEMux
    port map (
            O => \N__7941\,
            I => \N__7932\
        );

    \I__1774\ : Span4Mux_h
    port map (
            O => \N__7938\,
            I => \N__7928\
        );

    \I__1773\ : Span4Mux_h
    port map (
            O => \N__7935\,
            I => \N__7925\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__7932\,
            I => \N__7922\
        );

    \I__1771\ : CEMux
    port map (
            O => \N__7931\,
            I => \N__7919\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__7928\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1769\ : Odrv4
    port map (
            O => \N__7925\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__7922\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__7919\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\
        );

    \I__1766\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7907\,
            I => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\
        );

    \I__1764\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7901\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7901\,
            I => \N__7897\
        );

    \I__1762\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__1761\ : Span4Mux_h
    port map (
            O => \N__7897\,
            I => \N__7889\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7889\
        );

    \I__1759\ : Span4Mux_h
    port map (
            O => \N__7889\,
            I => \N__7886\
        );

    \I__1758\ : Sp12to4
    port map (
            O => \N__7886\,
            I => \N__7883\
        );

    \I__1757\ : Span12Mux_v
    port map (
            O => \N__7883\,
            I => \N__7880\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__7880\,
            I => \DRA_c_6\
        );

    \I__1755\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7874\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__7874\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7871\,
            I => \N__7868\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__7868\,
            I => \N__7865\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__7865\,
            I => \N__7861\
        );

    \I__1750\ : InMux
    port map (
            O => \N__7864\,
            I => \N__7858\
        );

    \I__1749\ : Span4Mux_h
    port map (
            O => \N__7861\,
            I => \N__7853\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__7858\,
            I => \N__7853\
        );

    \I__1747\ : Span4Mux_h
    port map (
            O => \N__7853\,
            I => \N__7850\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__7850\,
            I => \N__7847\
        );

    \I__1745\ : Span12Mux_v
    port map (
            O => \N__7847\,
            I => \N__7844\
        );

    \I__1744\ : Odrv12
    port map (
            O => \N__7844\,
            I => \DRA_c_5\
        );

    \I__1743\ : InMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__7838\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__7832\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1739\ : InMux
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7826\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__7820\,
            I => \N__7817\
        );

    \I__1735\ : Span4Mux_v
    port map (
            O => \N__7817\,
            I => \N__7813\
        );

    \I__1734\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__1733\ : Sp12to4
    port map (
            O => \N__7813\,
            I => \N__7805\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7810\,
            I => \N__7805\
        );

    \I__1731\ : Span12Mux_h
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1730\ : Span12Mux_v
    port map (
            O => \N__7802\,
            I => \N__7799\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__7799\,
            I => \DRA_c_1\
        );

    \I__1728\ : InMux
    port map (
            O => \N__7796\,
            I => \N__7793\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__7793\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1726\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7786\
        );

    \I__1725\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7783\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7783\,
            I => \N__7777\
        );

    \I__1722\ : Span4Mux_h
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__1721\ : Span12Mux_v
    port map (
            O => \N__7777\,
            I => \N__7771\
        );

    \I__1720\ : Sp12to4
    port map (
            O => \N__7774\,
            I => \N__7768\
        );

    \I__1719\ : Span12Mux_h
    port map (
            O => \N__7771\,
            I => \N__7765\
        );

    \I__1718\ : Span12Mux_v
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1717\ : Odrv12
    port map (
            O => \N__7765\,
            I => \DRA_c_2\
        );

    \I__1716\ : Odrv12
    port map (
            O => \N__7762\,
            I => \DRA_c_2\
        );

    \I__1715\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7754\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7754\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1713\ : InMux
    port map (
            O => \N__7751\,
            I => \N__7746\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7743\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7740\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7746\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__7743\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7740\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1707\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7729\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__7729\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__7726\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7721\,
            I => \N__7718\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__7718\,
            I => \N__7714\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__7714\,
            I => \N__7706\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7706\
        );

    \I__1698\ : Sp12to4
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1697\ : Span12Mux_v
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1696\ : Span12Mux_h
    port map (
            O => \N__7700\,
            I => \N__7697\
        );

    \I__1695\ : Odrv12
    port map (
            O => \N__7697\,
            I => \DRA_c_0\
        );

    \I__1694\ : CascadeMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__7682\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1689\ : IoInMux
    port map (
            O => \N__7679\,
            I => \N__7676\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__7676\,
            I => \N__7673\
        );

    \I__1687\ : Span4Mux_s3_v
    port map (
            O => \N__7673\,
            I => \N__7670\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__7670\,
            I => \N__7667\
        );

    \I__1685\ : Sp12to4
    port map (
            O => \N__7667\,
            I => \N__7664\
        );

    \I__1684\ : Odrv12
    port map (
            O => \N__7664\,
            I => \RASn_c\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7658\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__7655\,
            I => \N__7652\
        );

    \I__1680\ : Odrv4
    port map (
            O => \N__7652\,
            I => \U712_BYTE_ENABLE.un2_CLMBEnZ0\
        );

    \I__1679\ : IoInMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1677\ : Span4Mux_s3_h
    port map (
            O => \N__7643\,
            I => \N__7640\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1675\ : Sp12to4
    port map (
            O => \N__7637\,
            I => \N__7634\
        );

    \I__1674\ : Span12Mux_v
    port map (
            O => \N__7634\,
            I => \N__7631\
        );

    \I__1673\ : Odrv12
    port map (
            O => \N__7631\,
            I => \CLMBEn_c\
        );

    \I__1672\ : InMux
    port map (
            O => \N__7628\,
            I => \N__7623\
        );

    \I__1671\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7618\
        );

    \I__1670\ : InMux
    port map (
            O => \N__7626\,
            I => \N__7618\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7623\,
            I => \N__7613\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7618\,
            I => \N__7613\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__7613\,
            I => \N__7610\
        );

    \I__1666\ : Sp12to4
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1665\ : Span12Mux_h
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__1664\ : Span12Mux_v
    port map (
            O => \N__7604\,
            I => \N__7601\
        );

    \I__1663\ : Odrv12
    port map (
            O => \N__7601\,
            I => \CASUn_c\
        );

    \I__1662\ : IoInMux
    port map (
            O => \N__7598\,
            I => \N__7593\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__7597\,
            I => \N__7589\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__7596\,
            I => \N__7586\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7583\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7580\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7575\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7575\
        );

    \I__1655\ : Span12Mux_s5_v
    port map (
            O => \N__7583\,
            I => \N__7572\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7567\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7575\,
            I => \N__7567\
        );

    \I__1652\ : Span12Mux_v
    port map (
            O => \N__7572\,
            I => \N__7562\
        );

    \I__1651\ : Span4Mux_v
    port map (
            O => \N__7567\,
            I => \N__7559\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7566\,
            I => \N__7556\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7565\,
            I => \N__7553\
        );

    \I__1648\ : Odrv12
    port map (
            O => \N__7562\,
            I => \DBENn_c\
        );

    \I__1647\ : Odrv4
    port map (
            O => \N__7559\,
            I => \DBENn_c\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7556\,
            I => \DBENn_c\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7553\,
            I => \DBENn_c\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__7538\,
            I => \N__7535\
        );

    \I__1641\ : Odrv4
    port map (
            O => \N__7535\,
            I => \U712_BYTE_ENABLE.un2_CUUBEnZ0\
        );

    \I__1640\ : IoInMux
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__7529\,
            I => \N__7526\
        );

    \I__1638\ : IoSpan4Mux
    port map (
            O => \N__7526\,
            I => \N__7523\
        );

    \I__1637\ : IoSpan4Mux
    port map (
            O => \N__7523\,
            I => \N__7520\
        );

    \I__1636\ : Span4Mux_s3_h
    port map (
            O => \N__7520\,
            I => \N__7517\
        );

    \I__1635\ : Sp12to4
    port map (
            O => \N__7517\,
            I => \N__7514\
        );

    \I__1634\ : Odrv12
    port map (
            O => \N__7514\,
            I => \CUUBEn_c\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__7511\,
            I => \N__7508\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7504\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7507\,
            I => \N__7501\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7497\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7501\,
            I => \N__7494\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7500\,
            I => \N__7491\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__7497\,
            I => \N__7487\
        );

    \I__1626\ : Span12Mux_h
    port map (
            O => \N__7494\,
            I => \N__7482\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7491\,
            I => \N__7482\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7479\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__7487\,
            I => \REG_CYCLEm\
        );

    \I__1622\ : Odrv12
    port map (
            O => \N__7482\,
            I => \REG_CYCLEm\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7479\,
            I => \REG_CYCLEm\
        );

    \I__1620\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7466\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__7471\,
            I => \N__7462\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7470\,
            I => \N__7457\
        );

    \I__1617\ : InMux
    port map (
            O => \N__7469\,
            I => \N__7454\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7451\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7465\,
            I => \N__7444\
        );

    \I__1614\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7444\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7444\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__7460\,
            I => \N__7441\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__7457\,
            I => \N__7434\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7434\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__7451\,
            I => \N__7429\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7444\,
            I => \N__7429\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7426\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7440\,
            I => \N__7423\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7439\,
            I => \N__7420\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__7434\,
            I => \N__7417\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__7429\,
            I => \DMA_CYCLEm\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7426\,
            I => \DMA_CYCLEm\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__7423\,
            I => \DMA_CYCLEm\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7420\,
            I => \DMA_CYCLEm\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__7417\,
            I => \DMA_CYCLEm\
        );

    \I__1598\ : IoInMux
    port map (
            O => \N__7406\,
            I => \N__7403\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7403\,
            I => \N__7400\
        );

    \I__1596\ : Span4Mux_s2_v
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1595\ : Sp12to4
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1594\ : Span12Mux_s7_h
    port map (
            O => \N__7394\,
            I => \N__7391\
        );

    \I__1593\ : Span12Mux_v
    port map (
            O => \N__7391\,
            I => \N__7388\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__7388\,
            I => \N_52_i\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7385\,
            I => \N__7381\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7378\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7381\,
            I => \N__7375\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7378\,
            I => \N__7372\
        );

    \I__1587\ : Span4Mux_h
    port map (
            O => \N__7375\,
            I => \N__7369\
        );

    \I__1586\ : Sp12to4
    port map (
            O => \N__7372\,
            I => \N__7366\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__7369\,
            I => \N__7363\
        );

    \I__1584\ : Span12Mux_v
    port map (
            O => \N__7366\,
            I => \N__7358\
        );

    \I__1583\ : Sp12to4
    port map (
            O => \N__7363\,
            I => \N__7358\
        );

    \I__1582\ : Span12Mux_h
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__1581\ : Odrv12
    port map (
            O => \N__7355\,
            I => \DRA_c_7\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7349\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7343\,
            I => \U712_CHIP_RAM.N_37\
        );

    \I__1576\ : IoInMux
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7337\,
            I => \N__7334\
        );

    \I__1574\ : Span4Mux_s3_h
    port map (
            O => \N__7334\,
            I => \N__7331\
        );

    \I__1573\ : Span4Mux_v
    port map (
            O => \N__7331\,
            I => \N__7328\
        );

    \I__1572\ : Sp12to4
    port map (
            O => \N__7328\,
            I => \N__7325\
        );

    \I__1571\ : Span12Mux_h
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__1570\ : Odrv12
    port map (
            O => \N__7322\,
            I => \CMA_c_5\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7316\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7316\,
            I => \U712_CHIP_RAM.N_39\
        );

    \I__1567\ : IoInMux
    port map (
            O => \N__7313\,
            I => \N__7310\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__1565\ : IoSpan4Mux
    port map (
            O => \N__7307\,
            I => \N__7304\
        );

    \I__1564\ : Span4Mux_s2_h
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1563\ : Span4Mux_v
    port map (
            O => \N__7301\,
            I => \N__7298\
        );

    \I__1562\ : Sp12to4
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1561\ : Odrv12
    port map (
            O => \N__7295\,
            I => \CMA_c_7\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7289\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__1558\ : Span4Mux_v
    port map (
            O => \N__7286\,
            I => \N__7283\
        );

    \I__1557\ : Span4Mux_v
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1556\ : Sp12to4
    port map (
            O => \N__7280\,
            I => \N__7277\
        );

    \I__1555\ : Span12Mux_h
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1554\ : Odrv12
    port map (
            O => \N__7274\,
            I => \A_c_19\
        );

    \I__1553\ : IoInMux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1551\ : IoSpan4Mux
    port map (
            O => \N__7265\,
            I => \N__7262\
        );

    \I__1550\ : IoSpan4Mux
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1549\ : Span4Mux_s2_h
    port map (
            O => \N__7259\,
            I => \N__7256\
        );

    \I__1548\ : Sp12to4
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__7253\,
            I => \CMA_c_9\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__7244\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\
        );

    \I__1543\ : InMux
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7238\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7232\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_3\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1537\ : Span12Mux_v
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1536\ : Span12Mux_h
    port map (
            O => \N__7220\,
            I => \N__7217\
        );

    \I__1535\ : Odrv12
    port map (
            O => \N__7217\,
            I => \A_c_3\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7211\,
            I => \N__7208\
        );

    \I__1532\ : Span12Mux_v
    port map (
            O => \N__7208\,
            I => \N__7205\
        );

    \I__1531\ : Span12Mux_h
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__7202\,
            I => \A_c_10\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__7199\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7196\,
            I => \N__7193\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7193\,
            I => \N__7190\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__7190\,
            I => \U712_CHIP_RAM.N_33\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7184\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7184\,
            I => \N__7181\
        );

    \I__1523\ : Span4Mux_v
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__1522\ : Sp12to4
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__1521\ : Span12Mux_h
    port map (
            O => \N__7175\,
            I => \N__7172\
        );

    \I__1520\ : Odrv12
    port map (
            O => \N__7172\,
            I => \A_c_9\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7166\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7166\,
            I => \N__7163\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__7163\,
            I => \N__7160\
        );

    \I__1516\ : Sp12to4
    port map (
            O => \N__7160\,
            I => \N__7157\
        );

    \I__1515\ : Span12Mux_h
    port map (
            O => \N__7157\,
            I => \N__7154\
        );

    \I__1514\ : Span12Mux_v
    port map (
            O => \N__7154\,
            I => \N__7151\
        );

    \I__1513\ : Odrv12
    port map (
            O => \N__7151\,
            I => \A_c_2\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__7148\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1509\ : Odrv12
    port map (
            O => \N__7139\,
            I => \U712_CHIP_RAM.N_32\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7136\,
            I => \N__7129\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7135\,
            I => \N__7126\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__7134\,
            I => \N__7123\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7133\,
            I => \N__7120\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__7132\,
            I => \N__7117\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7129\,
            I => \N__7112\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7112\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7109\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7106\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7117\,
            I => \N__7103\
        );

    \I__1498\ : Span4Mux_h
    port map (
            O => \N__7112\,
            I => \N__7100\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7109\,
            I => \N__7095\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__7106\,
            I => \N__7095\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7103\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__7100\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1493\ : Odrv4
    port map (
            O => \N__7095\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1492\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1490\ : Odrv12
    port map (
            O => \N__7082\,
            I => \U712_BYTE_ENABLE.un2_CUMBEnZ0\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7079\,
            I => \N__7075\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7071\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7075\,
            I => \N__7068\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7065\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7071\,
            I => \N__7062\
        );

    \I__1484\ : Span4Mux_h
    port map (
            O => \N__7068\,
            I => \N__7057\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7065\,
            I => \N__7057\
        );

    \I__1482\ : Sp12to4
    port map (
            O => \N__7062\,
            I => \N__7054\
        );

    \I__1481\ : Sp12to4
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1480\ : Span12Mux_v
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1479\ : Span12Mux_h
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1478\ : Span12Mux_h
    port map (
            O => \N__7048\,
            I => \N__7040\
        );

    \I__1477\ : Span12Mux_v
    port map (
            O => \N__7045\,
            I => \N__7040\
        );

    \I__1476\ : Odrv12
    port map (
            O => \N__7040\,
            I => \CASLn_c\
        );

    \I__1475\ : IoInMux
    port map (
            O => \N__7037\,
            I => \N__7034\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1473\ : Span4Mux_s2_h
    port map (
            O => \N__7031\,
            I => \N__7028\
        );

    \I__1472\ : Sp12to4
    port map (
            O => \N__7028\,
            I => \N__7025\
        );

    \I__1471\ : Span12Mux_s5_v
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1470\ : Span12Mux_h
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__7019\,
            I => \CUMBEn_c\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7011\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7015\,
            I => \N__7008\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7014\,
            I => \N__7005\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7011\,
            I => \N__7000\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7008\,
            I => \N__7000\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7005\,
            I => \N__6996\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__7000\,
            I => \N__6993\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6990\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__6996\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\
        );

    \I__1459\ : Odrv4
    port map (
            O => \N__6993\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6990\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6978\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6973\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6981\,
            I => \N__6967\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6978\,
            I => \N__6964\
        );

    \I__1453\ : InMux
    port map (
            O => \N__6977\,
            I => \N__6961\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6958\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__6973\,
            I => \N__6955\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6972\,
            I => \N__6952\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6947\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6947\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6967\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6964\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6961\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6958\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__6955\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6952\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6947\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6929\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1438\ : Span12Mux_v
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1437\ : Span12Mux_h
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1436\ : Odrv12
    port map (
            O => \N__6920\,
            I => \A_c_16\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__6917\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1432\ : Span12Mux_v
    port map (
            O => \N__6908\,
            I => \N__6905\
        );

    \I__1431\ : Span12Mux_h
    port map (
            O => \N__6905\,
            I => \N__6902\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__6902\,
            I => \A_c_18\
        );

    \I__1429\ : IoInMux
    port map (
            O => \N__6899\,
            I => \N__6896\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__1427\ : Span4Mux_s2_v
    port map (
            O => \N__6893\,
            I => \N__6890\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1425\ : Span4Mux_v
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__1424\ : Odrv4
    port map (
            O => \N__6884\,
            I => \CMA_c_0\
        );

    \I__1423\ : IoInMux
    port map (
            O => \N__6881\,
            I => \N__6878\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1421\ : IoSpan4Mux
    port map (
            O => \N__6875\,
            I => \N__6872\
        );

    \I__1420\ : Span4Mux_s3_h
    port map (
            O => \N__6872\,
            I => \N__6869\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__6869\,
            I => \N__6866\
        );

    \I__1418\ : Span4Mux_v
    port map (
            O => \N__6866\,
            I => \N__6863\
        );

    \I__1417\ : Sp12to4
    port map (
            O => \N__6863\,
            I => \N__6860\
        );

    \I__1416\ : Odrv12
    port map (
            O => \N__6860\,
            I => \CMA_c_3\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6854\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1413\ : Span4Mux_h
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1412\ : Sp12to4
    port map (
            O => \N__6848\,
            I => \N__6845\
        );

    \I__1411\ : Span12Mux_v
    port map (
            O => \N__6845\,
            I => \N__6842\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__6842\,
            I => \N__6839\
        );

    \I__1409\ : Odrv12
    port map (
            O => \N__6839\,
            I => \A_c_5\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6827\
        );

    \I__1405\ : Span12Mux_v
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1404\ : Span12Mux_h
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1403\ : Odrv12
    port map (
            O => \N__6821\,
            I => \A_c_12\
        );

    \I__1402\ : InMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6815\,
            I => \U712_CHIP_RAM.N_35\
        );

    \I__1400\ : CascadeMux
    port map (
            O => \N__6812\,
            I => \N__6809\
        );

    \I__1399\ : InMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1397\ : Span4Mux_v
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1395\ : Sp12to4
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1394\ : Span12Mux_h
    port map (
            O => \N__6794\,
            I => \N__6791\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__6791\,
            I => \A_c_7\
        );

    \I__1392\ : InMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6785\,
            I => \N__6782\
        );

    \I__1390\ : Span12Mux_v
    port map (
            O => \N__6782\,
            I => \N__6779\
        );

    \I__1389\ : Span12Mux_h
    port map (
            O => \N__6779\,
            I => \N__6776\
        );

    \I__1388\ : Odrv12
    port map (
            O => \N__6776\,
            I => \A_c_14\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6770\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__6770\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_5\
        );

    \I__1385\ : CEMux
    port map (
            O => \N__6767\,
            I => \N__6764\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1383\ : Odrv12
    port map (
            O => \N__6761\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6758\,
            I => \N__6753\
        );

    \I__1381\ : InMux
    port map (
            O => \N__6757\,
            I => \N__6750\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6756\,
            I => \N__6747\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6753\,
            I => \N__6740\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6750\,
            I => \N__6740\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6747\,
            I => \N__6737\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6746\,
            I => \N__6731\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6731\
        );

    \I__1374\ : Span4Mux_v
    port map (
            O => \N__6740\,
            I => \N__6728\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__6737\,
            I => \N__6725\
        );

    \I__1372\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6722\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6731\,
            I => \N__6719\
        );

    \I__1370\ : Sp12to4
    port map (
            O => \N__6728\,
            I => \N__6712\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__6725\,
            I => \N__6712\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6722\,
            I => \N__6712\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__6719\,
            I => \N__6709\
        );

    \I__1366\ : Span12Mux_h
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__1364\ : Span12Mux_v
    port map (
            O => \N__6706\,
            I => \N__6700\
        );

    \I__1363\ : Odrv12
    port map (
            O => \N__6703\,
            I => \RnW_c\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__6700\,
            I => \RnW_c\
        );

    \I__1361\ : IoInMux
    port map (
            O => \N__6695\,
            I => \N__6692\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6692\,
            I => \N__6689\
        );

    \I__1359\ : Span4Mux_s3_v
    port map (
            O => \N__6689\,
            I => \N__6686\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__6686\,
            I => \N__6683\
        );

    \I__1357\ : Sp12to4
    port map (
            O => \N__6683\,
            I => \N__6679\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__6682\,
            I => \N__6675\
        );

    \I__1355\ : Span12Mux_s10_v
    port map (
            O => \N__6679\,
            I => \N__6672\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6669\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6666\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__6672\,
            I => \DBDIR_c\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6669\,
            I => \DBDIR_c\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6666\,
            I => \DBDIR_c\
        );

    \I__1349\ : IoInMux
    port map (
            O => \N__6659\,
            I => \N__6656\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6656\,
            I => \N__6653\
        );

    \I__1347\ : IoSpan4Mux
    port map (
            O => \N__6653\,
            I => \N__6650\
        );

    \I__1346\ : IoSpan4Mux
    port map (
            O => \N__6650\,
            I => \N__6647\
        );

    \I__1345\ : Span4Mux_s2_v
    port map (
            O => \N__6647\,
            I => \N__6644\
        );

    \I__1344\ : Sp12to4
    port map (
            O => \N__6644\,
            I => \N__6641\
        );

    \I__1343\ : Span12Mux_v
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1342\ : Odrv12
    port map (
            O => \N__6638\,
            I => \DRDDIR_0_i\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6621\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6618\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6609\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6609\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6609\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6609\
        );

    \I__1334\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6606\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6603\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6600\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6621\,
            I => \N__6591\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__6618\,
            I => \N__6591\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6609\,
            I => \N__6591\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6606\,
            I => \N__6591\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6588\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6584\
        );

    \I__1325\ : Span4Mux_v
    port map (
            O => \N__6591\,
            I => \N__6581\
        );

    \I__1324\ : Span4Mux_v
    port map (
            O => \N__6588\,
            I => \N__6578\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6587\,
            I => \N__6575\
        );

    \I__1322\ : Span12Mux_v
    port map (
            O => \N__6584\,
            I => \N__6570\
        );

    \I__1321\ : Sp12to4
    port map (
            O => \N__6581\,
            I => \N__6570\
        );

    \I__1320\ : Sp12to4
    port map (
            O => \N__6578\,
            I => \N__6565\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6575\,
            I => \N__6565\
        );

    \I__1318\ : Span12Mux_h
    port map (
            O => \N__6570\,
            I => \N__6562\
        );

    \I__1317\ : Span12Mux_h
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__1316\ : Odrv12
    port map (
            O => \N__6562\,
            I => \RESETn_c\
        );

    \I__1315\ : Odrv12
    port map (
            O => \N__6559\,
            I => \RESETn_c\
        );

    \I__1314\ : IoInMux
    port map (
            O => \N__6554\,
            I => \N__6551\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6548\
        );

    \I__1312\ : Span12Mux_s2_v
    port map (
            O => \N__6548\,
            I => \N__6545\
        );

    \I__1311\ : Odrv12
    port map (
            O => \N__6545\,
            I => \RESETn_c_i\
        );

    \I__1310\ : IoInMux
    port map (
            O => \N__6542\,
            I => \N__6539\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6539\,
            I => \N__6536\
        );

    \I__1308\ : Span4Mux_s0_v
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1307\ : Span4Mux_v
    port map (
            O => \N__6533\,
            I => \N__6530\
        );

    \I__1306\ : Span4Mux_v
    port map (
            O => \N__6530\,
            I => \N__6527\
        );

    \I__1305\ : Span4Mux_h
    port map (
            O => \N__6527\,
            I => \N__6524\
        );

    \I__1304\ : Odrv4
    port map (
            O => \N__6524\,
            I => \CRCSn_c\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6517\
        );

    \I__1302\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__6511\,
            I => \N__6502\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1297\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6497\
        );

    \I__1296\ : Span4Mux_h
    port map (
            O => \N__6502\,
            I => \N__6494\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6489\
        );

    \I__1294\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6489\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6497\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1292\ : Odrv4
    port map (
            O => \N__6494\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__6489\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__6482\,
            I => \N__6479\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6476\
        );

    \I__1288\ : IoSpan4Mux
    port map (
            O => \N__6476\,
            I => \N__6473\
        );

    \I__1287\ : Sp12to4
    port map (
            O => \N__6473\,
            I => \N__6470\
        );

    \I__1286\ : Span12Mux_s9_v
    port map (
            O => \N__6470\,
            I => \N__6467\
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__6467\,
            I => \CMA_c_10\
        );

    \I__1284\ : IoInMux
    port map (
            O => \N__6464\,
            I => \N__6461\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6461\,
            I => \N__6458\
        );

    \I__1282\ : Span4Mux_s2_v
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1281\ : Span4Mux_v
    port map (
            O => \N__6455\,
            I => \N__6452\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__6452\,
            I => \N__6449\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__6449\,
            I => \CMA_c_1\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6443\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6443\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6437\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6437\,
            I => \N__6433\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1273\ : Span4Mux_v
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1271\ : Sp12to4
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1270\ : Sp12to4
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__1269\ : Span12Mux_h
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1268\ : Span12Mux_v
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1267\ : Span12Mux_v
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1266\ : Span12Mux_h
    port map (
            O => \N__6412\,
            I => \N__6406\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__6409\,
            I => \DRA_c_3\
        );

    \I__1264\ : Odrv12
    port map (
            O => \N__6406\,
            I => \DRA_c_3\
        );

    \I__1263\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6398\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__6395\,
            I => \U712_CHIP_RAM.N_47_cascade_\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1259\ : LocalMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__6386\,
            I => \U712_CHIP_RAM.N_89\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6379\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6376\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6379\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6376\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__6368\,
            I => \U712_CHIP_RAM.N_100\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__6365\,
            I => \U712_CHIP_RAM.N_100_cascade_\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6362\,
            I => \N__6358\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6358\,
            I => \U712_CHIP_RAM.N_101\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.N_101\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6340\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6343\,
            I => \N__6337\
        );

    \I__1242\ : Span4Mux_v
    port map (
            O => \N__6340\,
            I => \N__6334\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__1239\ : Span4Mux_v
    port map (
            O => \N__6331\,
            I => \N__6325\
        );

    \I__1238\ : Sp12to4
    port map (
            O => \N__6328\,
            I => \N__6320\
        );

    \I__1237\ : Sp12to4
    port map (
            O => \N__6325\,
            I => \N__6320\
        );

    \I__1236\ : Span12Mux_h
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1235\ : Odrv12
    port map (
            O => \N__6317\,
            I => \AWEn_c\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6308\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__6305\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6298\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__6298\,
            I => \N__6292\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6295\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__6292\,
            I => \U712_CHIP_RAM.WRITE_CYCLEZ0\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6284\,
            I => \N__6279\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__6283\,
            I => \N__6276\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6265\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6279\,
            I => \N__6262\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6259\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6256\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6274\,
            I => \N__6249\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6249\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6272\,
            I => \N__6249\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6271\,
            I => \N__6246\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6243\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6238\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6238\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6265\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1210\ : Odrv12
    port map (
            O => \N__6262\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6259\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__6256\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6249\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6246\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6243\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6238\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__6221\,
            I => \N__6217\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6211\
        );

    \I__1200\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6208\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__6211\,
            I => \N__6205\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6194\
        );

    \I__1197\ : Span4Mux_v
    port map (
            O => \N__6205\,
            I => \N__6191\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6204\,
            I => \N__6188\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6185\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6182\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6179\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6176\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6173\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6168\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6168\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__6194\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__6191\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6188\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6185\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6182\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__6179\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6173\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6168\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6144\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6140\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__6147\,
            I => \N__6137\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6134\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6128\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6125\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6122\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__6134\,
            I => \N__6119\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6133\,
            I => \N__6114\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6114\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6131\,
            I => \N__6111\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6128\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6125\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6122\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__6119\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.N_56\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__6098\,
            I => \N__6094\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6090\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6087\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6082\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6079\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6087\,
            I => \N__6076\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6071\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6085\,
            I => \N__6071\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6082\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6079\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6076\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6071\,
            I => \U712_CHIP_RAM.N_42\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__6062\,
            I => \N__6053\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6046\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6046\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6035\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6030\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6030\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6056\,
            I => \N__6027\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6024\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6052\,
            I => \N__6019\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6019\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6016\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6011\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6011\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6006\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6042\,
            I => \N__6006\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6003\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6040\,
            I => \N__5996\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6039\,
            I => \N__5996\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6038\,
            I => \N__5996\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__5991\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__6030\,
            I => \N__5991\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6027\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__6024\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__6019\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1126\ : Odrv4
    port map (
            O => \N__6016\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6011\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6006\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6003\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__5996\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1121\ : Odrv4
    port map (
            O => \N__5991\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__5972\,
            I => \N__5959\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5953\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5953\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5946\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5946\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5940\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5933\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5933\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5933\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5929\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5924\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5924\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5958\,
            I => \N__5921\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5953\,
            I => \N__5918\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5913\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5913\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5946\,
            I => \N__5910\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5907\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5902\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5902\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5897\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5897\
        );

    \I__1098\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5894\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5929\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5924\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__5921\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1094\ : Odrv4
    port map (
            O => \N__5918\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5913\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__5910\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5907\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1090\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1089\ : Odrv4
    port map (
            O => \N__5897\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5894\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__5873\,
            I => \U712_CHIP_RAM.N_42_cascade_\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5863\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5856\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__5863\,
            I => \N__5853\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5850\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5843\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5860\,
            I => \N__5843\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5859\,
            I => \N__5843\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__5856\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__5853\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5850\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5843\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__5831\,
            I => \N__5828\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__5828\,
            I => \N__5824\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__1070\ : Odrv4
    port map (
            O => \N__5824\,
            I => \U712_CHIP_RAM.N_98\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5821\,
            I => \U712_CHIP_RAM.N_98\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5813\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5813\,
            I => \N__5810\
        );

    \I__1066\ : Span12Mux_v
    port map (
            O => \N__5810\,
            I => \N__5807\
        );

    \I__1065\ : Span12Mux_h
    port map (
            O => \N__5807\,
            I => \N__5804\
        );

    \I__1064\ : Odrv12
    port map (
            O => \N__5804\,
            I => \A_c_15\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__5801\,
            I => \N__5798\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5798\,
            I => \N__5795\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5792\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__5792\,
            I => \N__5789\
        );

    \I__1059\ : Span4Mux_v
    port map (
            O => \N__5789\,
            I => \N__5786\
        );

    \I__1058\ : Sp12to4
    port map (
            O => \N__5786\,
            I => \N__5783\
        );

    \I__1057\ : Span12Mux_h
    port map (
            O => \N__5783\,
            I => \N__5780\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__5780\,
            I => \A_c_8\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5774\,
            I => \U712_CHIP_RAM.N_38\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5768\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__5768\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_6\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5759\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5752\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5749\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5746\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5759\,
            I => \N__5743\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5740\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5737\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5732\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5732\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5752\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__5749\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5746\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1039\ : Odrv4
    port map (
            O => \N__5743\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__5740\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5732\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5710\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__1032\ : Span4Mux_v
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5707\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__5704\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__1027\ : Span4Mux_h
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__5690\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5681\,
            I => \N__5677\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__1021\ : Span4Mux_h
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5674\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__5671\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1018\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5663\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__1016\ : Span4Mux_h
    port map (
            O => \N__5660\,
            I => \N__5657\
        );

    \I__1015\ : Odrv4
    port map (
            O => \N__5657\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__1014\ : InMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5651\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__5648\,
            I => \N__5645\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5645\,
            I => \N__5641\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5638\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5641\,
            I => \N__5635\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\
        );

    \I__1007\ : Odrv4
    port map (
            O => \N__5635\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5626\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5629\,
            I => \N__5623\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5623\,
            I => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5618\,
            I => \N__5613\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5608\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5616\,
            I => \N__5608\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5613\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5608\,
            I => \U712_CHIP_RAM.REFRESH_CYCLEZ0\
        );

    \I__997\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5599\
        );

    \I__996\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5599\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5596\,
            I => \U712_CHIP_RAM.N_47\
        );

    \I__993\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5588\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\
        );

    \I__991\ : InMux
    port map (
            O => \N__5585\,
            I => \N__5580\
        );

    \I__990\ : InMux
    port map (
            O => \N__5584\,
            I => \N__5575\
        );

    \I__989\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5575\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5580\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5575\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__5570\,
            I => \N__5566\
        );

    \I__985\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__984\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5563\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5560\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__981\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5548\
        );

    \I__979\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__5548\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5545\,
            I => \U712_CHIP_RAM.N_57\
        );

    \I__976\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5537\,
            I => \U712_BYTE_ENABLE.un2_CLLBEnZ0\
        );

    \I__974\ : IoInMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__972\ : IoSpan4Mux
    port map (
            O => \N__5528\,
            I => \N__5525\
        );

    \I__971\ : Span4Mux_s2_v
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__970\ : Sp12to4
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__969\ : Span12Mux_v
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__5516\,
            I => \CLLBEn_c\
        );

    \I__967\ : InMux
    port map (
            O => \N__5513\,
            I => \N__5510\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5510\,
            I => \U712_CHIP_RAM.DMA_CYCLE_7\
        );

    \I__965\ : InMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5504\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0\
        );

    \I__963\ : IoInMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__961\ : IoSpan4Mux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__960\ : IoSpan4Mux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__958\ : Span12Mux_s9_h
    port map (
            O => \N__5486\,
            I => \N__5483\
        );

    \I__957\ : Odrv12
    port map (
            O => \N__5483\,
            I => \CMA_c_6\
        );

    \I__956\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5477\,
            I => \N__5474\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__5474\,
            I => \U712_CHIP_RAM.un1_CMA31_0_i\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__5471\,
            I => \U712_CHIP_RAM.N_44_cascade_\
        );

    \I__952\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5463\
        );

    \I__951\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5460\
        );

    \I__950\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5457\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5463\,
            I => \U712_CHIP_RAM.N_93\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__5460\,
            I => \U712_CHIP_RAM.N_93\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5457\,
            I => \U712_CHIP_RAM.N_93\
        );

    \I__946\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5446\
        );

    \I__945\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5443\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5446\,
            I => \U712_CHIP_RAM.N_13\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5443\,
            I => \U712_CHIP_RAM.N_13\
        );

    \I__942\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5435\,
            I => \U712_CHIP_RAM.N_65\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__5432\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5426\,
            I => \U712_CHIP_RAM.N_62\
        );

    \I__937\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5417\
        );

    \I__936\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5414\
        );

    \I__935\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5409\
        );

    \I__934\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5409\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5417\,
            I => \N__5402\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5402\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5409\,
            I => \N__5402\
        );

    \I__930\ : Odrv4
    port map (
            O => \N__5402\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\
        );

    \I__929\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5394\
        );

    \I__928\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5389\
        );

    \I__927\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5389\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5394\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__5389\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__923\ : InMux
    port map (
            O => \N__5381\,
            I => \N__5375\
        );

    \I__922\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5368\
        );

    \I__921\ : InMux
    port map (
            O => \N__5379\,
            I => \N__5368\
        );

    \I__920\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5368\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5375\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5368\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__5363\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\
        );

    \I__916\ : InMux
    port map (
            O => \N__5360\,
            I => \N__5350\
        );

    \I__915\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5350\
        );

    \I__914\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5350\
        );

    \I__913\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5347\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5347\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\
        );

    \I__910\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5339\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5339\,
            I => \U712_CHIP_RAM.N_75\
        );

    \I__908\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5332\
        );

    \I__907\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5329\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5332\,
            I => \U712_CHIP_RAM.N_60\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5329\,
            I => \U712_CHIP_RAM.N_60\
        );

    \I__904\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5321\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5321\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1\
        );

    \I__902\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5315\,
            I => \U712_CHIP_RAM.N_77\
        );

    \I__900\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__5309\,
            I => \U712_CHIP_RAM.N_40\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__5306\,
            I => \U712_CHIP_RAM.N_62_cascade_\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__5303\,
            I => \U712_CHIP_RAM.N_13_cascade_\
        );

    \I__896\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__893\ : Sp12to4
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__892\ : Span12Mux_h
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__891\ : Span12Mux_v
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__890\ : Odrv12
    port map (
            O => \N__5282\,
            I => \A_c_4\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__888\ : InMux
    port map (
            O => \N__5276\,
            I => \N__5273\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__884\ : Span12Mux_h
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__5261\,
            I => \A_c_11\
        );

    \I__882\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5255\,
            I => \U712_CHIP_RAM.N_34\
        );

    \I__880\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5249\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__878\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5243\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_2\
        );

    \I__876\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5237\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__874\ : SRMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__872\ : Odrv4
    port map (
            O => \N__5228\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__5225\,
            I => \U712_CHIP_RAM.N_74_cascade_\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__5222\,
            I => \U712_CHIP_RAM.N_50_cascade_\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5219\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\
        );

    \I__868\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5213\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5213\,
            I => \U712_CHIP_RAM.N_58\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__5210\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_\
        );

    \I__865\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5204\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5200\
        );

    \I__863\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5197\
        );

    \I__862\ : Span12Mux_h
    port map (
            O => \N__5200\,
            I => \N__5192\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5192\
        );

    \I__860\ : Span12Mux_h
    port map (
            O => \N__5192\,
            I => \N__5189\
        );

    \I__859\ : Span12Mux_v
    port map (
            O => \N__5189\,
            I => \N__5186\
        );

    \I__858\ : Odrv12
    port map (
            O => \N__5186\,
            I => \SIZ_c_1\
        );

    \I__857\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5173\
        );

    \I__856\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5173\
        );

    \I__855\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5173\
        );

    \I__854\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5170\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5173\,
            I => \N__5165\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5165\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__5165\,
            I => \N__5161\
        );

    \I__850\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5158\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__5158\,
            I => \N__5152\
        );

    \I__847\ : Sp12to4
    port map (
            O => \N__5155\,
            I => \N__5147\
        );

    \I__846\ : Span12Mux_v
    port map (
            O => \N__5152\,
            I => \N__5147\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__5147\,
            I => \A_c_0\
        );

    \I__844\ : InMux
    port map (
            O => \N__5144\,
            I => \N__5141\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__5141\,
            I => \U712_BYTE_ENABLE.LLBE_0_0_tz\
        );

    \I__842\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5132\
        );

    \I__841\ : InMux
    port map (
            O => \N__5137\,
            I => \N__5125\
        );

    \I__840\ : InMux
    port map (
            O => \N__5136\,
            I => \N__5125\
        );

    \I__839\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5125\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5132\,
            I => \U712_BYTE_ENABLE.LW_TRANS_0\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5125\,
            I => \U712_BYTE_ENABLE.LW_TRANS_0\
        );

    \I__836\ : CascadeMux
    port map (
            O => \N__5120\,
            I => \U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_\
        );

    \I__835\ : CascadeMux
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__834\ : InMux
    port map (
            O => \N__5114\,
            I => \N__5110\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__5113\,
            I => \N__5106\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5102\
        );

    \I__831\ : InMux
    port map (
            O => \N__5109\,
            I => \N__5095\
        );

    \I__830\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5095\
        );

    \I__829\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5095\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__5102\,
            I => \N__5090\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5095\,
            I => \N__5090\
        );

    \I__826\ : Span4Mux_v
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__825\ : Span4Mux_v
    port map (
            O => \N__5087\,
            I => \N__5084\
        );

    \I__824\ : Sp12to4
    port map (
            O => \N__5084\,
            I => \N__5081\
        );

    \I__823\ : Span12Mux_h
    port map (
            O => \N__5081\,
            I => \N__5078\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__5078\,
            I => \A_c_1\
        );

    \I__821\ : IoInMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5072\,
            I => \N__5069\
        );

    \I__819\ : Odrv12
    port map (
            O => \N__5069\,
            I => \CMA_c_2\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \U712_CHIP_RAM.N_58_cascade_\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__5063\,
            I => \U712_CHIP_RAM.N_40_cascade_\
        );

    \I__816\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5057\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.N_99_cascade_\
        );

    \I__813\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5048\,
            I => \U712_CHIP_RAM.N_85\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__5045\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_\
        );

    \I__810\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5039\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__5036\,
            I => \U712_CHIP_RAM.N_65_cascade_\
        );

    \I__807\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5030\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5027\,
            I => \U712_CHIP_RAM.N_49_cascade_\
        );

    \I__804\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5020\
        );

    \I__803\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5017\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5020\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5017\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__800\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5008\
        );

    \I__799\ : InMux
    port map (
            O => \N__5011\,
            I => \N__5005\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5008\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5005\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__5000\,
            I => \N__4996\
        );

    \I__795\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4993\
        );

    \I__794\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4990\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4993\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4990\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__791\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4981\
        );

    \I__790\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4978\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4981\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__4978\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__787\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4969\
        );

    \I__786\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4969\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4966\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__783\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4957\
        );

    \I__782\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4954\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4957\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4954\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__779\ : CascadeMux
    port map (
            O => \N__4949\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_\
        );

    \I__778\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4943\,
            I => \N__4939\
        );

    \I__776\ : IoInMux
    port map (
            O => \N__4942\,
            I => \N__4936\
        );

    \I__775\ : Span12Mux_h
    port map (
            O => \N__4939\,
            I => \N__4933\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__4936\,
            I => \N__4930\
        );

    \I__773\ : Span12Mux_v
    port map (
            O => \N__4933\,
            I => \N__4927\
        );

    \I__772\ : IoSpan4Mux
    port map (
            O => \N__4930\,
            I => \N__4924\
        );

    \I__771\ : Odrv12
    port map (
            O => \N__4927\,
            I => \RAMENn_c\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__4924\,
            I => \RAMENn_c\
        );

    \I__769\ : CascadeMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__768\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4913\,
            I => \N__4909\
        );

    \I__766\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4906\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__4909\,
            I => \N__4900\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4906\,
            I => \N__4900\
        );

    \I__763\ : InMux
    port map (
            O => \N__4905\,
            I => \N__4897\
        );

    \I__762\ : Span4Mux_v
    port map (
            O => \N__4900\,
            I => \N__4894\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4891\
        );

    \I__760\ : Sp12to4
    port map (
            O => \N__4894\,
            I => \N__4888\
        );

    \I__759\ : Span12Mux_h
    port map (
            O => \N__4891\,
            I => \N__4885\
        );

    \I__758\ : Span12Mux_h
    port map (
            O => \N__4888\,
            I => \N__4882\
        );

    \I__757\ : Span12Mux_v
    port map (
            O => \N__4885\,
            I => \N__4879\
        );

    \I__756\ : Span12Mux_v
    port map (
            O => \N__4882\,
            I => \N__4876\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__4879\,
            I => \TSn_c\
        );

    \I__754\ : Odrv12
    port map (
            O => \N__4876\,
            I => \TSn_c\
        );

    \I__753\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4867\
        );

    \I__752\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4863\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4867\,
            I => \N__4860\
        );

    \I__750\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4857\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4863\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__4860\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4857\,
            I => \U712_REG_SM_DBR_SYNC_1\
        );

    \I__746\ : CascadeMux
    port map (
            O => \N__4850\,
            I => \N__4846\
        );

    \I__745\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4840\
        );

    \I__744\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4840\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__4845\,
            I => \N__4836\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4840\,
            I => \N__4833\
        );

    \I__741\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4830\
        );

    \I__740\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4827\
        );

    \I__739\ : Odrv12
    port map (
            O => \N__4833\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4830\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__4827\,
            I => \U712_REG_SM_DBR_SYNC_0\
        );

    \I__736\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4814\
        );

    \I__735\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4814\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__733\ : CascadeMux
    port map (
            O => \N__4811\,
            I => \U712_CHIP_RAM.N_57_cascade_\
        );

    \I__732\ : InMux
    port map (
            O => \N__4808\,
            I => \bfn_10_7_0_\
        );

    \I__731\ : InMux
    port map (
            O => \N__4805\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__730\ : InMux
    port map (
            O => \N__4802\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__729\ : InMux
    port map (
            O => \N__4799\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__728\ : InMux
    port map (
            O => \N__4796\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__727\ : InMux
    port map (
            O => \N__4793\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__726\ : InMux
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__725\ : InMux
    port map (
            O => \N__4787\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__724\ : ClkMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__723\ : GlobalMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__722\ : gio2CtrlBuf
    port map (
            O => \N__4778\,
            I => \C1_c_g\
        );

    \I__721\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4772\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__718\ : Sp12to4
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__717\ : Span12Mux_h
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__716\ : Span12Mux_v
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__715\ : Odrv12
    port map (
            O => \N__4757\,
            I => \DBRn_c\
        );

    \I__714\ : InMux
    port map (
            O => \N__4754\,
            I => \N__4749\
        );

    \I__713\ : InMux
    port map (
            O => \N__4753\,
            I => \N__4746\
        );

    \I__712\ : InMux
    port map (
            O => \N__4752\,
            I => \N__4743\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4749\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4746\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4743\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__708\ : CascadeMux
    port map (
            O => \N__4736\,
            I => \N__4731\
        );

    \I__707\ : InMux
    port map (
            O => \N__4735\,
            I => \N__4728\
        );

    \I__706\ : InMux
    port map (
            O => \N__4734\,
            I => \N__4723\
        );

    \I__705\ : InMux
    port map (
            O => \N__4731\,
            I => \N__4723\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4728\,
            I => \N__4720\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4723\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__702\ : Odrv4
    port map (
            O => \N__4720\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__701\ : CEMux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4712\,
            I => \N__4709\
        );

    \I__699\ : Span4Mux_h
    port map (
            O => \N__4709\,
            I => \N__4706\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__4706\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_0\
        );

    \I__697\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4700\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4700\,
            I => \U712_REG_SM.LDS_OUT_2_0_0\
        );

    \I__695\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4694\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4690\
        );

    \I__693\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4686\
        );

    \I__692\ : Span4Mux_h
    port map (
            O => \N__4690\,
            I => \N__4683\
        );

    \I__691\ : InMux
    port map (
            O => \N__4689\,
            I => \N__4680\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4686\,
            I => \N__4677\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__4683\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__4680\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__4677\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__686\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4666\
        );

    \I__685\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4663\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4666\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4663\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__682\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4655\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__4652\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \N__4645\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__4648\,
            I => \N__4641\
        );

    \I__677\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4638\
        );

    \I__676\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4635\
        );

    \I__675\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4632\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4638\,
            I => \N__4629\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__4635\,
            I => \N__4624\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4632\,
            I => \N__4624\
        );

    \I__671\ : Sp12to4
    port map (
            O => \N__4629\,
            I => \N__4621\
        );

    \I__670\ : Span12Mux_h
    port map (
            O => \N__4624\,
            I => \N__4618\
        );

    \I__669\ : Span12Mux_v
    port map (
            O => \N__4621\,
            I => \N__4615\
        );

    \I__668\ : Span12Mux_v
    port map (
            O => \N__4618\,
            I => \N__4612\
        );

    \I__667\ : Odrv12
    port map (
            O => \N__4615\,
            I => \SIZ_c_0\
        );

    \I__666\ : Odrv12
    port map (
            O => \N__4612\,
            I => \SIZ_c_0\
        );

    \I__665\ : InMux
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__663\ : Odrv4
    port map (
            O => \N__4601\,
            I => \TACK_EN_i_ess\
        );

    \I__662\ : IoInMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__660\ : Span4Mux_s0_h
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__659\ : Sp12to4
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__658\ : Span12Mux_v
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__656\ : Odrv12
    port map (
            O => \N__4580\,
            I => \N_614_i\
        );

    \I__655\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4574\,
            I => \U712_CHIP_RAM.N_36\
        );

    \I__653\ : IoInMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__651\ : Span4Mux_s3_h
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__650\ : Span4Mux_v
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__647\ : Sp12to4
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__646\ : Odrv12
    port map (
            O => \N__4550\,
            I => \CMA_c_4\
        );

    \I__645\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4544\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__643\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4537\
        );

    \I__642\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4534\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4537\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4534\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_1\
        );

    \I__639\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4526\,
            I => \U712_REG_SM.N_188\
        );

    \I__637\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4519\
        );

    \I__636\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4519\,
            I => \N__4511\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__4516\,
            I => \N__4511\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__4511\,
            I => \REG_TACK\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__4505\,
            I => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\
        );

    \I__630\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4495\
        );

    \I__628\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__4495\,
            I => \N__4487\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4492\,
            I => \N__4487\
        );

    \I__625\ : Span4Mux_v
    port map (
            O => \N__4487\,
            I => \N__4484\
        );

    \I__624\ : Sp12to4
    port map (
            O => \N__4484\,
            I => \N__4481\
        );

    \I__623\ : Span12Mux_h
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__622\ : Odrv12
    port map (
            O => \N__4478\,
            I => \REGSPACEn_c\
        );

    \I__621\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4471\
        );

    \I__620\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4468\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4471\,
            I => \N__4464\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__4468\,
            I => \N__4461\
        );

    \I__617\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4458\
        );

    \I__616\ : Odrv4
    port map (
            O => \N__4464\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__4461\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4458\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1\
        );

    \I__613\ : CascadeMux
    port map (
            O => \N__4451\,
            I => \N__4446\
        );

    \I__612\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4443\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__4449\,
            I => \N__4440\
        );

    \I__610\ : InMux
    port map (
            O => \N__4446\,
            I => \N__4437\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4443\,
            I => \N__4434\
        );

    \I__608\ : InMux
    port map (
            O => \N__4440\,
            I => \N__4431\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4437\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__606\ : Odrv4
    port map (
            O => \N__4434\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4431\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_0\
        );

    \I__604\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4420\
        );

    \I__603\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4417\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__4420\,
            I => \CPU_TACKm\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4417\,
            I => \CPU_TACKm\
        );

    \I__600\ : CascadeMux
    port map (
            O => \N__4412\,
            I => \N__4406\
        );

    \I__599\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4403\
        );

    \I__598\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4400\
        );

    \I__597\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4395\
        );

    \I__596\ : InMux
    port map (
            O => \N__4406\,
            I => \N__4395\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4403\,
            I => \N__4392\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4389\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4395\,
            I => \N__4386\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__4392\,
            I => \N__4383\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__4389\,
            I => \N__4378\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__4386\,
            I => \N__4378\
        );

    \I__589\ : Sp12to4
    port map (
            O => \N__4383\,
            I => \N__4375\
        );

    \I__588\ : Span4Mux_h
    port map (
            O => \N__4378\,
            I => \N__4372\
        );

    \I__587\ : Span12Mux_h
    port map (
            O => \N__4375\,
            I => \N__4367\
        );

    \I__586\ : Sp12to4
    port map (
            O => \N__4372\,
            I => \N__4367\
        );

    \I__585\ : Span12Mux_v
    port map (
            O => \N__4367\,
            I => \N__4364\
        );

    \I__584\ : Odrv12
    port map (
            O => \N__4364\,
            I => \CLK40_OUT_i\
        );

    \I__583\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4355\
        );

    \I__582\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4355\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4350\
        );

    \I__580\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4345\
        );

    \I__579\ : InMux
    port map (
            O => \N__4353\,
            I => \N__4345\
        );

    \I__578\ : Odrv4
    port map (
            O => \N__4350\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4345\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__576\ : CascadeMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__575\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4333\
        );

    \I__574\ : InMux
    port map (
            O => \N__4336\,
            I => \N__4330\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4333\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4330\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__571\ : InMux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__569\ : Odrv4
    port map (
            O => \N__4319\,
            I => \U712_REG_SM.UDS_OUT_2_0_0\
        );

    \I__568\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4312\
        );

    \I__567\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4309\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4312\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4309\,
            I => \U712_REG_SM.LDS_OUTZ0\
        );

    \I__564\ : IoInMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__562\ : IoSpan4Mux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__561\ : IoSpan4Mux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__560\ : Span4Mux_s2_v
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__559\ : Sp12to4
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__558\ : Span12Mux_v
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__557\ : Odrv12
    port map (
            O => \N__4283\,
            I => \U712_REG_SM_un1_LDSn_i\
        );

    \I__556\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4277\,
            I => \N__4273\
        );

    \I__554\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4270\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__4273\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4270\,
            I => \U712_REG_SM.UDS_OUTZ0\
        );

    \I__551\ : InMux
    port map (
            O => \N__4265\,
            I => \N__4261\
        );

    \I__550\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4258\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4261\,
            I => \N__4252\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__547\ : InMux
    port map (
            O => \N__4257\,
            I => \N__4249\
        );

    \I__546\ : Odrv12
    port map (
            O => \N__4252\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4249\,
            I => \U712_REG_SM.DS_ENZ0\
        );

    \I__544\ : IoInMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__542\ : IoSpan4Mux
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__541\ : IoSpan4Mux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__539\ : Span12Mux_v
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__4226\,
            I => \U712_REG_SM_un1_UDSn_i\
        );

    \I__537\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__535\ : Span4Mux_v
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__534\ : Sp12to4
    port map (
            O => \N__4214\,
            I => \N__4211\
        );

    \I__533\ : Odrv12
    port map (
            O => \N__4211\,
            I => \A_c_13\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__4208\,
            I => \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\
        );

    \I__531\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4202\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__529\ : Span4Mux_h
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__4196\,
            I => \N__4193\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__4190\,
            I => \A_c_6\
        );

    \I__525\ : InMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4184\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__4181\,
            I => \N__4175\
        );

    \I__522\ : InMux
    port map (
            O => \N__4180\,
            I => \N__4172\
        );

    \I__521\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4169\
        );

    \I__520\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4166\
        );

    \I__519\ : InMux
    port map (
            O => \N__4175\,
            I => \N__4163\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4172\,
            I => \N__4160\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4169\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4163\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__514\ : Odrv4
    port map (
            O => \N__4160\,
            I => \U712_REG_SM.N_163_0\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__4151\,
            I => \N__4147\
        );

    \I__512\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4144\
        );

    \I__511\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4141\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4135\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4141\,
            I => \N__4129\
        );

    \I__508\ : InMux
    port map (
            O => \N__4140\,
            I => \N__4126\
        );

    \I__507\ : InMux
    port map (
            O => \N__4139\,
            I => \N__4121\
        );

    \I__506\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4121\
        );

    \I__505\ : Span4Mux_h
    port map (
            O => \N__4135\,
            I => \N__4118\
        );

    \I__504\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4111\
        );

    \I__503\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4111\
        );

    \I__502\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4111\
        );

    \I__501\ : Odrv4
    port map (
            O => \N__4129\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4126\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__4121\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__4118\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4111\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__496\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4097\,
            I => \U712_REG_SM.N_186\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4094\,
            I => \U712_REG_SM.N_176_0_cascade_\
        );

    \I__493\ : InMux
    port map (
            O => \N__4091\,
            I => \N__4085\
        );

    \I__492\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4080\
        );

    \I__491\ : InMux
    port map (
            O => \N__4089\,
            I => \N__4080\
        );

    \I__490\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4077\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4085\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4080\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4077\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__486\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4063\
        );

    \I__485\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__484\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4060\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4063\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4060\,
            I => \U712_REG_SM.C3_SYNCZ0Z_2\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__480\ : InMux
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__4049\,
            I => \N__4045\
        );

    \I__478\ : InMux
    port map (
            O => \N__4048\,
            I => \N__4042\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__4045\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4042\,
            I => \U712_REG_SM.N_157_0\
        );

    \I__475\ : InMux
    port map (
            O => \N__4037\,
            I => \N__4029\
        );

    \I__474\ : InMux
    port map (
            O => \N__4036\,
            I => \N__4024\
        );

    \I__473\ : InMux
    port map (
            O => \N__4035\,
            I => \N__4024\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4034\,
            I => \N__4021\
        );

    \I__471\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4017\
        );

    \I__470\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4014\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__4029\,
            I => \N__4009\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4024\,
            I => \N__4009\
        );

    \I__467\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4006\
        );

    \I__466\ : InMux
    port map (
            O => \N__4020\,
            I => \N__4003\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4017\,
            I => \N__4000\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__4014\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__4009\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4006\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4003\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__4000\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__459\ : CascadeMux
    port map (
            O => \N__3989\,
            I => \N__3982\
        );

    \I__458\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3979\
        );

    \I__457\ : InMux
    port map (
            O => \N__3987\,
            I => \N__3976\
        );

    \I__456\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3973\
        );

    \I__455\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3968\
        );

    \I__454\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3968\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3979\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3976\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3973\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3968\,
            I => \U712_REG_SM.C1_SYNCZ0Z_2\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__3959\,
            I => \U712_REG_SM.N_157_0_cascade_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__447\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3945\
        );

    \I__446\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3942\
        );

    \I__445\ : InMux
    port map (
            O => \N__3951\,
            I => \N__3939\
        );

    \I__444\ : InMux
    port map (
            O => \N__3950\,
            I => \N__3932\
        );

    \I__443\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3932\
        );

    \I__442\ : InMux
    port map (
            O => \N__3948\,
            I => \N__3932\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__3945\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3942\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3939\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3932\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__437\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3920\,
            I => \U712_REG_SM.N_176_0\
        );

    \I__435\ : CascadeMux
    port map (
            O => \N__3917\,
            I => \N__3912\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__3916\,
            I => \N__3909\
        );

    \I__433\ : InMux
    port map (
            O => \N__3915\,
            I => \N__3906\
        );

    \I__432\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3901\
        );

    \I__431\ : InMux
    port map (
            O => \N__3909\,
            I => \N__3901\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3906\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3901\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__428\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3893\,
            I => \N__3887\
        );

    \I__426\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3880\
        );

    \I__425\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3880\
        );

    \I__424\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3880\
        );

    \I__423\ : Odrv4
    port map (
            O => \N__3887\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3880\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_5\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__3875\,
            I => \N__3871\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__3874\,
            I => \N__3868\
        );

    \I__419\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3865\
        );

    \I__418\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3861\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3865\,
            I => \N__3858\
        );

    \I__416\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3855\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3861\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__414\ : Odrv4
    port map (
            O => \N__3858\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3855\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__412\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3845\,
            I => \U712_REG_SM.N_192\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__408\ : Span4Mux_s0_h
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__407\ : Span4Mux_h
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__406\ : Sp12to4
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__405\ : Span12Mux_v
    port map (
            O => \N__3827\,
            I => \N__3823\
        );

    \I__404\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3820\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__3823\,
            I => \TACK_OUTn\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3820\,
            I => \TACK_OUTn\
        );

    \I__401\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3811\
        );

    \I__400\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3807\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3811\,
            I => \N__3803\
        );

    \I__398\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3800\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3807\,
            I => \N__3797\
        );

    \I__396\ : InMux
    port map (
            O => \N__3806\,
            I => \N__3794\
        );

    \I__395\ : Odrv12
    port map (
            O => \N__3803\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3800\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__393\ : Odrv4
    port map (
            O => \N__3797\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3794\,
            I => \U712_REG_SM.N_171_0\
        );

    \I__391\ : IoInMux
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__389\ : Span12Mux_s4_v
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__388\ : Odrv12
    port map (
            O => \N__3776\,
            I => \VBENn_c\
        );

    \I__387\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3766\
        );

    \I__385\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3763\
        );

    \I__384\ : Odrv4
    port map (
            O => \N__3766\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3763\,
            I => \U712_REG_SM.N_162_0\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__3758\,
            I => \U712_REG_SM.N_171_0_cascade_\
        );

    \I__381\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3752\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3752\,
            I => \U712_REG_SM.RnW_m\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__3749\,
            I => \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__3746\,
            I => \N__3742\
        );

    \I__377\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3738\
        );

    \I__376\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3735\
        );

    \I__375\ : InMux
    port map (
            O => \N__3741\,
            I => \N__3732\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3738\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3735\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3732\,
            I => \U712_REG_SM.N_165_0\
        );

    \I__371\ : CascadeMux
    port map (
            O => \N__3725\,
            I => \U712_REG_SM.N_167_0_cascade_\
        );

    \I__370\ : InMux
    port map (
            O => \N__3722\,
            I => \N__3713\
        );

    \I__369\ : InMux
    port map (
            O => \N__3721\,
            I => \N__3713\
        );

    \I__368\ : InMux
    port map (
            O => \N__3720\,
            I => \N__3713\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3713\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_2\
        );

    \I__366\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3704\
        );

    \I__365\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3704\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3704\,
            I => \U712_REG_SM.N_167_0\
        );

    \I__363\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3696\
        );

    \I__362\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3693\
        );

    \I__361\ : InMux
    port map (
            O => \N__3699\,
            I => \N__3690\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3696\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__3693\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3690\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_6\
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__3683\,
            I => \U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_\
        );

    \I__356\ : InMux
    port map (
            O => \N__3680\,
            I => \N__3677\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3677\,
            I => \N__3673\
        );

    \I__354\ : IoInMux
    port map (
            O => \N__3676\,
            I => \N__3670\
        );

    \I__353\ : Span4Mux_v
    port map (
            O => \N__3673\,
            I => \N__3667\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3670\,
            I => \N__3664\
        );

    \I__351\ : Sp12to4
    port map (
            O => \N__3667\,
            I => \N__3661\
        );

    \I__350\ : Span4Mux_s3_h
    port map (
            O => \N__3664\,
            I => \N__3658\
        );

    \I__349\ : Span12Mux_h
    port map (
            O => \N__3661\,
            I => \N__3653\
        );

    \I__348\ : Sp12to4
    port map (
            O => \N__3658\,
            I => \N__3653\
        );

    \I__347\ : Span12Mux_v
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3650\,
            I => \C1_c\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__3647\,
            I => \U712_REG_SM.N_162_0_cascade_\
        );

    \I__344\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3641\,
            I => \N__3636\
        );

    \I__342\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3631\
        );

    \I__341\ : InMux
    port map (
            O => \N__3639\,
            I => \N__3631\
        );

    \I__340\ : Odrv4
    port map (
            O => \N__3636\,
            I => \U712_REG_SM.N_166_0\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3631\,
            I => \U712_REG_SM.N_166_0\
        );

    \I__338\ : InMux
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3623\,
            I => \N__3620\
        );

    \I__336\ : Span12Mux_h
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__335\ : Span12Mux_v
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__334\ : Odrv12
    port map (
            O => \N__3614\,
            I => \C3_c\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__3611\,
            I => \U712_REG_SM.REG_TACK_7_0_cascade_\
        );

    \I__332\ : InMux
    port map (
            O => \N__3608\,
            I => \N__3604\
        );

    \I__331\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3601\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__3604\,
            I => \U712_REG_SM.un1_STATE_COUNT_5_0_1\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3601\,
            I => \U712_REG_SM.un1_STATE_COUNT_5_0_1\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__3596\,
            I => \U712_REG_SM.N_183_cascade_\
        );

    \I__327\ : IoInMux
    port map (
            O => \N__3593\,
            I => \N__3590\
        );

    \I__326\ : LocalMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__325\ : Odrv12
    port map (
            O => \N__3587\,
            I => \CLK40_OUT_i_i\
        );

    \I__324\ : IoInMux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__322\ : Span4Mux_s2_v
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__321\ : Span4Mux_v
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__320\ : Span4Mux_h
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__319\ : Odrv4
    port map (
            O => \N__3569\,
            I => \CLK80_OUT_i_i\
        );

    \I__318\ : IoInMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__317\ : LocalMux
    port map (
            O => \N__3563\,
            I => \N__3559\
        );

    \I__316\ : IoInMux
    port map (
            O => \N__3562\,
            I => \N__3556\
        );

    \I__315\ : IoSpan4Mux
    port map (
            O => \N__3559\,
            I => \N__3553\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3556\,
            I => \N__3550\
        );

    \I__313\ : Sp12to4
    port map (
            O => \N__3553\,
            I => \N__3547\
        );

    \I__312\ : IoSpan4Mux
    port map (
            O => \N__3550\,
            I => \N__3544\
        );

    \I__311\ : Span12Mux_s6_v
    port map (
            O => \N__3547\,
            I => \N__3541\
        );

    \I__310\ : Sp12to4
    port map (
            O => \N__3544\,
            I => \N__3538\
        );

    \I__309\ : Span12Mux_v
    port map (
            O => \N__3541\,
            I => \N__3535\
        );

    \I__308\ : Span12Mux_s6_v
    port map (
            O => \N__3538\,
            I => \N__3532\
        );

    \I__307\ : Span12Mux_h
    port map (
            O => \N__3535\,
            I => \N__3526\
        );

    \I__306\ : Span12Mux_v
    port map (
            O => \N__3532\,
            I => \N__3526\
        );

    \I__305\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3523\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__3526\,
            I => \ASn_c\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__3523\,
            I => \ASn_c\
        );

    \I__302\ : IoInMux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__3515\,
            I => \N__3512\
        );

    \I__300\ : IoSpan4Mux
    port map (
            O => \N__3512\,
            I => \N__3509\
        );

    \I__299\ : Span4Mux_s2_v
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__298\ : Sp12to4
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__297\ : Span12Mux_v
    port map (
            O => \N__3503\,
            I => \N__3500\
        );

    \I__296\ : Odrv12
    port map (
            O => \N__3500\,
            I => \CLK40_IN_c\
        );

    \IN_MUX_bfv_10_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_7_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__6554\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3676\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLK40C_obuf_RNO_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4411\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9287\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_OUT_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__3810\,
            in1 => \N__3531\,
            in2 => \_gnd_net_\,
            in3 => \N__4474\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9270\,
            ce => 'H',
            sr => \N__9064\
        );

    \U712_REG_SM.STATE_COUNT_5_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3607\,
            in2 => \_gnd_net_\,
            in3 => \N__3644\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9270\,
            ce => 'H',
            sr => \N__9064\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__3891\,
            in1 => \N__6746\,
            in2 => \N__3917\,
            in3 => \N__3639\,
            lcout => OPEN,
            ltout => \U712_REG_SM.REG_TACK_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000001111"
        )
    port map (
            in0 => \N__4523\,
            in1 => \N__3701\,
            in2 => \N__3611\,
            in3 => \N__3608\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9274\,
            ce => 'H',
            sr => \N__9058\
        );

    \U712_REG_SM.STATE_COUNT_RNIFFKI2_4_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__3890\,
            in1 => \N__4139\,
            in2 => \N__3916\,
            in3 => \N__4178\,
            lcout => \U712_REG_SM.un1_STATE_COUNT_5_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_6_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4037\,
            in1 => \N__3745\,
            in2 => \N__3956\,
            in3 => \N__3988\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_6_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000001100"
        )
    port map (
            in0 => \N__3892\,
            in1 => \N__3700\,
            in2 => \N__3596\,
            in3 => \N__3640\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9274\,
            ce => 'H',
            sr => \N__9058\
        );

    \U712_REG_SM.DS_EN_RNO_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6745\,
            in2 => \_gnd_net_\,
            in3 => \N__4138\,
            lcout => \U712_REG_SM.RnW_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIQU741_2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4089\,
            in1 => \N__4069\,
            in2 => \_gnd_net_\,
            in3 => \N__4133\,
            lcout => \U712_REG_SM.N_165_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9278\,
            ce => 'H',
            sr => \N__9051\
        );

    \U712_REG_SM.C1_SYNC_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3950\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9278\,
            ce => 'H',
            sr => \N__9051\
        );

    \U712_REG_SM.STATE_COUNT_RNI81E81_6_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__3949\,
            in1 => \N__3699\,
            in2 => \N__4034\,
            in3 => \N__3985\,
            lcout => OPEN,
            ltout => \U712_REG_SM.DS_EN_0_sqmuxa_1_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI20MC2_6_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3683\,
            in3 => \N__3741\,
            lcout => \U712_REG_SM.DS_EN_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3680\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9278\,
            ce => 'H',
            sr => \N__9051\
        );

    \U712_REG_SM.C1_SYNC_RNI9DCD1_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4033\,
            in1 => \N__4132\,
            in2 => \N__3989\,
            in3 => \N__3948\,
            lcout => \U712_REG_SM.N_162_0\,
            ltout => \U712_REG_SM.N_162_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIIDN62_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__4070\,
            in1 => \_gnd_net_\,
            in2 => \N__3647\,
            in3 => \N__4090\,
            lcout => \U712_REG_SM.N_166_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_2_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4091\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9281\,
            ce => 'H',
            sr => \N__9041\
        );

    \U712_REG_SM.C3_SYNC_0_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__3626\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9281\,
            ce => 'H',
            sr => \N__9041\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4032\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9281\,
            ce => 'H',
            sr => \N__9041\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4670\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9283\,
            ce => 'H',
            sr => \N__9033\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7500\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8861\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__4529\,
            in1 => \N__3773\,
            in2 => \N__4055\,
            in3 => \N__4450\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9265\,
            ce => 'H',
            sr => \N__9059\
        );

    \U712_REG_SM.STATE_COUNT_RNITQLC2_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4540\,
            in1 => \N__3769\,
            in2 => \_gnd_net_\,
            in3 => \N__4048\,
            lcout => \U712_REG_SM.N_171_0\,
            ltout => \U712_REG_SM.N_171_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_RNO_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__3720\,
            in1 => \N__3709\,
            in2 => \N__3758\,
            in3 => \N__4467\,
            lcout => OPEN,
            ltout => \U712_REG_SM.un1_LDS_OUT_0_sqmuxa_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DS_EN_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__3755\,
            in1 => \N__4036\,
            in2 => \N__3749\,
            in3 => \N__4257\,
            lcout => \U712_REG_SM.DS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9271\,
            ce => 'H',
            sr => \N__9052\
        );

    \U712_REG_SM.C1_SYNC_RNIIDN62_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4035\,
            in1 => \N__3987\,
            in2 => \N__3746\,
            in3 => \N__3952\,
            lcout => \U712_REG_SM.N_167_0\,
            ltout => \U712_REG_SM.N_167_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3721\,
            in2 => \N__3725\,
            in3 => \N__3806\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9271\,
            ce => 'H',
            sr => \N__9052\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011011000"
        )
    port map (
            in0 => \N__3722\,
            in1 => \N__3710\,
            in2 => \N__3874\,
            in3 => \N__4100\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9271\,
            ce => 'H',
            sr => \N__9052\
        );

    \U712_REG_SM.STATE_COUNT_RNIVAPS2_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__4839\,
            in2 => \N__4181\,
            in3 => \N__3864\,
            lcout => \U712_REG_SM.N_176_0\,
            ltout => \U712_REG_SM.N_176_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4094\,
            in3 => \N__4140\,
            lcout => \U712_REG_SM.N_192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI90BP_2_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4088\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4068\,
            lcout => \U712_REG_SM.N_157_0\,
            ltout => \U712_REG_SM.N_157_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI1FQR1_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4020\,
            in1 => \N__3986\,
            in2 => \N__3959\,
            in3 => \N__3951\,
            lcout => \U712_REG_SM.N_163_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111000100"
        )
    port map (
            in0 => \N__4179\,
            in1 => \N__3923\,
            in2 => \N__4151\,
            in3 => \N__3915\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9275\,
            ce => 'H',
            sr => \N__9042\
        );

    \U712_REG_SM.REG_CYCLE_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011100100"
        )
    port map (
            in0 => \N__3896\,
            in1 => \N__7490\,
            in2 => \N__3875\,
            in3 => \N__3848\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9279\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_REG_SM.UDS_OUT_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__4325\,
            in1 => \N__4276\,
            in2 => \N__4649\,
            in3 => \N__3814\,
            lcout => \U712_REG_SM.UDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9279\,
            ce => 'H',
            sr => \N__9034\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111000100"
        )
    port map (
            in0 => \N__4361\,
            in1 => \N__3826\,
            in2 => \N__4412\,
            in3 => \N__4689\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9282\,
            ce => 'H',
            sr => \N__9022\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4409\,
            in2 => \_gnd_net_\,
            in3 => \N__4360\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9282\,
            ce => 'H',
            sr => \N__9022\
        );

    \U712_REG_SM.LDS_OUT_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__4703\,
            in1 => \N__4315\,
            in2 => \N__4648\,
            in3 => \N__3815\,
            lcout => \U712_REG_SM.LDS_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9282\,
            ce => 'H',
            sr => \N__9022\
        );

    \U712_REG_SM.UDS_OUT_RNO_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6736\,
            in2 => \_gnd_net_\,
            in3 => \N__5164\,
            lcout => \U712_REG_SM.UDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDS_OUT_RNIL31J_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4316\,
            lcout => \U712_REG_SM_un1_LDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDS_OUT_RNIUP9B_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4280\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4265\,
            lcout => \U712_REG_SM_un1_UDSn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__4187\,
            in1 => \N__8856\,
            in2 => \N__8133\,
            in3 => \N__4547\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8857\,
            in1 => \N__4223\,
            in2 => \N__4208\,
            in3 => \N__4205\,
            lcout => \U712_CHIP_RAM.N_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_5_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7871\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9252\,
            ce => \N__8285\,
            sr => \N__9060\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4180\,
            in1 => \N__4870\,
            in2 => \N__4850\,
            in3 => \N__4150\,
            lcout => \U712_REG_SM.N_186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4849\,
            lcout => \U712_REG_SM_DBR_SYNC_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9259\,
            ce => 'H',
            sr => \N__9053\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101111"
        )
    port map (
            in0 => \N__4905\,
            in1 => \N__4498\,
            in2 => \N__4449\,
            in3 => \N__4541\,
            lcout => \U712_REG_SM.N_188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN6_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4522\,
            in2 => \_gnd_net_\,
            in3 => \N__4423\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => \U712_CYCLE_TERM.TACK_EN6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6625\,
            in1 => \N__4752\,
            in2 => \N__4508\,
            in3 => \N__4336\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_45_0_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__9119\,
            in1 => \_gnd_net_\,
            in2 => \N__4505\,
            in3 => \_gnd_net_\,
            lcout => \U712_CYCLE_TERM.N_45_0_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011111000"
        )
    port map (
            in0 => \N__4658\,
            in1 => \N__4734\,
            in2 => \N__4340\,
            in3 => \N__4353\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__4912\,
            in1 => \N__4502\,
            in2 => \N__4451\,
            in3 => \N__4475\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__4424\,
            in1 => \N__5033\,
            in2 => \N__6221\,
            in3 => \N__8864\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010001100"
        )
    port map (
            in0 => \N__4354\,
            in1 => \N__4753\,
            in2 => \N__4736\,
            in3 => \N__4410\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4697\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CHIP_RAM.DBR_SYNC_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4775\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM_DBR_SYNC_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9272\,
            ce => 'H',
            sr => \N__9035\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__6587\,
            in1 => \N__4754\,
            in2 => \_gnd_net_\,
            in3 => \N__4735\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9276\,
            ce => \N__4715\,
            sr => \N__9023\
        );

    \U712_REG_SM.LDS_OUT_RNO_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6756\,
            lcout => \U712_REG_SM.LDS_OUT_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4693\,
            in2 => \_gnd_net_\,
            in3 => \N__4669\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_a3_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LW_TRANS_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__5203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4644\,
            lcout => \U712_BYTE_ENABLE.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_obuft_RNO_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4607\,
            lcout => \N_614_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8433\,
            in1 => \N__4577\,
            in2 => \_gnd_net_\,
            in3 => \N__8552\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9236\,
            ce => \N__8646\,
            sr => \N__9065\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7789\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9245\,
            ce => \N__7961\,
            sr => \N__9061\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8330\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9245\,
            ce => \N__7961\,
            sr => \N__9061\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4985\,
            in2 => \_gnd_net_\,
            in3 => \N__4808\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_10_7_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5012\,
            in2 => \_gnd_net_\,
            in3 => \N__4805\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5024\,
            in2 => \_gnd_net_\,
            in3 => \N__4802\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5713\,
            in2 => \_gnd_net_\,
            in3 => \N__4799\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4999\,
            in2 => \_gnd_net_\,
            in3 => \N__4796\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4961\,
            in2 => \_gnd_net_\,
            in3 => \N__4793\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4973\,
            in2 => \_gnd_net_\,
            in3 => \N__4790\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5680\,
            in2 => \_gnd_net_\,
            in3 => \N__4787\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4784\,
            ce => 'H',
            sr => \N__5234\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000100000"
        )
    port map (
            in0 => \N__5966\,
            in1 => \N__5763\,
            in2 => \N__6635\,
            in3 => \N__5335\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_49_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__5357\,
            in1 => \_gnd_net_\,
            in2 => \N__5027\,
            in3 => \N__6507\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9253\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__5023\,
            in1 => \N__5011\,
            in2 => \N__5000\,
            in3 => \N__4984\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4972\,
            in2 => \_gnd_net_\,
            in3 => \N__4960\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_2_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__6058\,
            in2 => \_gnd_net_\,
            in3 => \N__6203\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISSMN4_3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001000"
        )
    port map (
            in0 => \N__6149\,
            in1 => \N__5467\,
            in2 => \N__4949\,
            in3 => \N__6275\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_0_2_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6057\,
            in1 => \N__5964\,
            in2 => \_gnd_net_\,
            in3 => \N__6202\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101011"
        )
    port map (
            in0 => \N__4820\,
            in1 => \N__4946\,
            in2 => \N__4919\,
            in3 => \N__8848\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9260\,
            ce => 'H',
            sr => \N__9036\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI17BM1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__4866\,
            in1 => \N__7133\,
            in2 => \N__4845\,
            in3 => \N__4819\,
            lcout => \U712_CHIP_RAM.N_57\,
            ltout => \U712_CHIP_RAM.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0V852_2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4811\,
            in3 => \N__6199\,
            lcout => \U712_CHIP_RAM.N_58\,
            ltout => \U712_CHIP_RAM.N_58_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSC34_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5952\,
            in1 => \N__6044\,
            in2 => \N__5066\,
            in3 => \N__5466\,
            lcout => \U712_CHIP_RAM.N_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIN7BL3_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000010"
        )
    port map (
            in0 => \N__6382\,
            in1 => \N__5951\,
            in2 => \N__5870\,
            in3 => \N__6392\,
            lcout => \U712_CHIP_RAM.N_40\,
            ltout => \U712_CHIP_RAM.N_40_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUB006_0_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6045\,
            in2 => \N__5063\,
            in3 => \N__6143\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_99_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3F0BF_0_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__6631\,
            in1 => \N__5060\,
            in2 => \N__5054\,
            in3 => \N__5051\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__5756\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6039\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQ4PC1_1_2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6040\,
            in1 => \N__5958\,
            in2 => \_gnd_net_\,
            in3 => \N__6204\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_3_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6133\,
            in1 => \N__5758\,
            in2 => \N__5045\,
            in3 => \N__6273\,
            lcout => \U712_CHIP_RAM.N_65\,
            ltout => \U712_CHIP_RAM.N_65_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__5944\,
            in1 => \N__5042\,
            in2 => \N__5036\,
            in3 => \N__6097\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_5_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__5422\,
            in1 => \N__5399\,
            in2 => \N__5384\,
            in3 => \N__6274\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__9116\,
            in1 => \_gnd_net_\,
            in2 => \N__5219\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITJ7E1_0_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5755\,
            in1 => \N__6038\,
            in2 => \_gnd_net_\,
            in3 => \N__5943\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_a2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI7Q5U5_3_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6272\,
            in1 => \N__5216\,
            in2 => \N__5210\,
            in3 => \N__6132\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CUMBEn_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000000"
        )
    port map (
            in0 => \N__5144\,
            in1 => \N__5138\,
            in2 => \N__5117\,
            in3 => \N__8850\,
            lcout => \U712_BYTE_ENABLE.un2_CUMBEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CLMBEn_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010100000000"
        )
    port map (
            in0 => \N__5136\,
            in1 => \N__5182\,
            in2 => \N__5113\,
            in3 => \N__8852\,
            lcout => \U712_BYTE_ENABLE.un2_CLMBEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CUUBEn_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__5183\,
            in1 => \N__5137\,
            in2 => \N__8863\,
            in3 => \N__5109\,
            lcout => \U712_BYTE_ENABLE.un2_CUUBEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_0_tz_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5181\,
            lcout => \U712_BYTE_ENABLE.LLBE_0_0_tz\,
            ltout => \U712_BYTE_ENABLE.LLBE_0_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un2_CLLBEn_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000100010"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__5135\,
            in2 => \N__5120\,
            in3 => \N__5105\,
            lcout => \U712_BYTE_ENABLE.un2_CLLBEnZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8556\,
            in1 => \N__5258\,
            in2 => \_gnd_net_\,
            in3 => \N__8442\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9231\,
            ce => \N__8645\,
            sr => \N__9069\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__5300\,
            in1 => \N__8862\,
            in2 => \N__5279\,
            in3 => \N__5246\,
            lcout => \U712_CHIP_RAM.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__5240\,
            in1 => \N__8826\,
            in2 => \N__8118\,
            in3 => \N__5252\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_3_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6440\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9237\,
            ce => \N__8281\,
            sr => \N__9054\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000010011"
        )
    port map (
            in0 => \N__8510\,
            in1 => \N__6501\,
            in2 => \N__8061\,
            in3 => \N__8389\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6500\,
            in1 => \N__8509\,
            in2 => \N__8417\,
            in3 => \N__8025\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6628\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5834\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_74_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__5359\,
            in1 => \N__5342\,
            in2 => \N__5225\,
            in3 => \N__8416\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__6629\,
            in1 => \N__5318\,
            in2 => \N__5648\,
            in3 => \N__6362\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_50_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111100000101"
        )
    port map (
            in0 => \N__5358\,
            in1 => \_gnd_net_\,
            in2 => \N__5222\,
            in3 => \N__8060\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6059\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111110101"
        )
    port map (
            in0 => \N__5360\,
            in1 => \N__5336\,
            in2 => \N__8557\,
            in3 => \N__6627\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9249\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5967\,
            in1 => \N__6302\,
            in2 => \_gnd_net_\,
            in3 => \N__5468\,
            lcout => \U712_CHIP_RAM.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVGRT_2_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6201\,
            in2 => \_gnd_net_\,
            in3 => \N__6270\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_1_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI264TB_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__6361\,
            in1 => \N__5827\,
            in2 => \_gnd_net_\,
            in3 => \N__6970\,
            lcout => \U712_CHIP_RAM.N_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5602\,
            in1 => \N__5324\,
            in2 => \N__5972\,
            in3 => \N__6093\,
            lcout => \U712_CHIP_RAM.N_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIKLSF6_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__6051\,
            in1 => \N__5312\,
            in2 => \N__6148\,
            in3 => \N__9117\,
            lcout => \U712_CHIP_RAM.N_62\,
            ltout => \U712_CHIP_RAM.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI13TLG_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__6971\,
            in1 => \N__5762\,
            in2 => \N__5306\,
            in3 => \N__7015\,
            lcout => \U712_CHIP_RAM.N_13\,
            ltout => \U712_CHIP_RAM.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__5423\,
            in1 => \_gnd_net_\,
            in2 => \N__5303\,
            in3 => \N__6282\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001000110000"
        )
    port map (
            in0 => \N__5962\,
            in1 => \N__5449\,
            in2 => \N__6220\,
            in3 => \N__6052\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9254\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__5862\,
            in1 => \N__5630\,
            in2 => \_gnd_net_\,
            in3 => \N__5618\,
            lcout => \U712_CHIP_RAM.N_44\,
            ltout => \U712_CHIP_RAM.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNIOG801_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__6626\,
            in1 => \_gnd_net_\,
            in2 => \N__5471\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__6056\,
            in1 => \N__5963\,
            in2 => \_gnd_net_\,
            in3 => \N__5450\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000001"
        )
    port map (
            in0 => \N__5764\,
            in1 => \N__5551\,
            in2 => \N__6062\,
            in3 => \N__6976\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__5438\,
            in1 => \_gnd_net_\,
            in2 => \N__5432\,
            in3 => \N__5429\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__5397\,
            in2 => \N__5570\,
            in3 => \N__5378\,
            lcout => \U712_CHIP_RAM.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001101010"
        )
    port map (
            in0 => \N__5380\,
            in1 => \N__5421\,
            in2 => \N__6287\,
            in3 => \N__9111\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIIP2_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5420\,
            in1 => \N__5398\,
            in2 => \N__6283\,
            in3 => \N__5379\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER_13_c6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9112\,
            in2 => \N__5363\,
            in3 => \N__5584\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__5591\,
            in1 => \N__5585\,
            in2 => \N__9122\,
            in3 => \N__5569\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9261\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9110\,
            in2 => \_gnd_net_\,
            in3 => \N__6999\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBDIR_RNO_0_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5555\,
            in2 => \_gnd_net_\,
            in3 => \N__5765\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101010101"
        )
    port map (
            in0 => \N__5540\,
            in1 => \N__7079\,
            in2 => \N__7460\,
            in3 => \N__7566\,
            lcout => \CLLBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIH4474_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7135\,
            in2 => \_gnd_net_\,
            in3 => \N__6972\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__7014\,
            in1 => \N__7565\,
            in2 => \N__7694\,
            in3 => \N__5513\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9273\,
            ce => 'H',
            sr => \N__9013\
        );

    \U712_CHIP_RAM.DBDIR_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011000111110000"
        )
    port map (
            in0 => \N__6982\,
            in1 => \N__6343\,
            in2 => \N__6682\,
            in3 => \N__5507\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9273\,
            ce => 'H',
            sr => \N__9013\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__5777\,
            in1 => \N__8575\,
            in2 => \_gnd_net_\,
            in3 => \N__8454\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9230\,
            ce => \N__8616\,
            sr => \N__9057\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9120\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5480\,
            lcout => \U712_CHIP_RAM.un1_CMA31_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000110011"
        )
    port map (
            in0 => \N__5816\,
            in1 => \N__5771\,
            in2 => \N__5801\,
            in3 => \N__8838\,
            lcout => \U712_CHIP_RAM.N_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8787\,
            in1 => \N__6446\,
            in2 => \N__8114\,
            in3 => \N__6401\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6060\,
            in1 => \N__5757\,
            in2 => \_gnd_net_\,
            in3 => \N__5970\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_1_sqmuxa_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6JQ74_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000001"
        )
    port map (
            in0 => \N__6061\,
            in1 => \N__5603\,
            in2 => \N__6098\,
            in3 => \N__5971\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__5717\,
            in1 => \N__5699\,
            in2 => \N__5687\,
            in3 => \N__5666\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => 'H',
            sr => \N__9018\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__8794\,
            in1 => \N__5654\,
            in2 => \_gnd_net_\,
            in3 => \N__7470\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => 'H',
            sr => \N__9018\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__5617\,
            in1 => \N__5644\,
            in2 => \_gnd_net_\,
            in3 => \N__6983\,
            lcout => \U712_CHIP_RAM.REFRESH_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => 'H',
            sr => \N__9018\
        );

    \U712_CHIP_RAM.REFRESH_CYCLE_START_RNI27CG_0_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5859\,
            in1 => \N__5629\,
            in2 => \_gnd_net_\,
            in3 => \N__5616\,
            lcout => \U712_CHIP_RAM.N_47\,
            ltout => \U712_CHIP_RAM.N_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVE5T1_2_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6197\,
            in1 => \N__5932\,
            in2 => \N__6395\,
            in3 => \N__6268\,
            lcout => \U712_CHIP_RAM.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5861\,
            in1 => \N__6371\,
            in2 => \_gnd_net_\,
            in3 => \N__6383\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9248\,
            ce => 'H',
            sr => \N__9018\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI0CV43_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5945\,
            in1 => \N__6041\,
            in2 => \N__6147\,
            in3 => \N__5860\,
            lcout => \U712_CHIP_RAM.N_100\,
            ltout => \U712_CHIP_RAM.N_100_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVSQ24_2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100000"
        )
    port map (
            in0 => \N__6269\,
            in1 => \_gnd_net_\,
            in2 => \N__6365\,
            in3 => \N__6198\,
            lcout => \U712_CHIP_RAM.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__7439\,
            in1 => \N__6758\,
            in2 => \N__6350\,
            in3 => \N__8849\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001001110"
        )
    port map (
            in0 => \N__6314\,
            in1 => \N__6301\,
            in2 => \N__6305\,
            in3 => \N__6086\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9251\,
            ce => 'H',
            sr => \N__9014\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6042\,
            in1 => \N__5968\,
            in2 => \_gnd_net_\,
            in3 => \N__6085\,
            lcout => \U712_CHIP_RAM.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9VIP2_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6271\,
            in1 => \N__6200\,
            in2 => \_gnd_net_\,
            in3 => \N__6131\,
            lcout => \U712_CHIP_RAM.N_42\,
            ltout => \U712_CHIP_RAM.N_42_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000101"
        )
    port map (
            in0 => \N__6043\,
            in1 => \N__5969\,
            in2 => \N__5873\,
            in3 => \N__5866\,
            lcout => \U712_CHIP_RAM.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7136\,
            in2 => \_gnd_net_\,
            in3 => \N__6977\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9258\,
            ce => \N__6767\,
            sr => \N__9012\
        );

    \U712_BUFFERS.DRDDIR_0_i_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__6757\,
            in1 => \N__6678\,
            in2 => \N__7511\,
            in3 => \N__7440\,
            lcout => \DRDDIR_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6624\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6520\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9232\,
            ce => 'H',
            sr => \N__9070\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_13_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8574\,
            in1 => \N__8119\,
            in2 => \N__8471\,
            in3 => \N__6521\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9233\,
            ce => \N__8621\,
            sr => \N__9066\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100000001"
        )
    port map (
            in0 => \N__8123\,
            in1 => \N__8576\,
            in2 => \N__8472\,
            in3 => \N__7196\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9234\,
            ce => \N__8617\,
            sr => \N__9062\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_7_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7385\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9238\,
            ce => \N__8280\,
            sr => \N__9055\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9246\,
            ce => \N__7957\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7904\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9246\,
            ce => \N__7957\,
            sr => \N__9043\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__7016\,
            in1 => \N__8768\,
            in2 => \N__7132\,
            in3 => \N__6981\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9255\,
            ce => 'H',
            sr => \N__9024\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7250\,
            in1 => \N__8841\,
            in2 => \N__8134\,
            in3 => \N__7352\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001101"
        )
    port map (
            in0 => \N__8842\,
            in1 => \N__6932\,
            in2 => \N__6917\,
            in3 => \N__6914\,
            lcout => \U712_CHIP_RAM.N_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8583\,
            in1 => \N__7145\,
            in2 => \_gnd_net_\,
            in3 => \N__8461\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => \N__8653\,
            sr => \N__9067\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8584\,
            in1 => \N__6818\,
            in2 => \_gnd_net_\,
            in3 => \N__8462\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9239\,
            ce => \N__8653\,
            sr => \N__9067\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110011"
        )
    port map (
            in0 => \N__6857\,
            in1 => \N__8844\,
            in2 => \N__6836\,
            in3 => \N__7235\,
            lcout => \U712_CHIP_RAM.N_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010110010001"
        )
    port map (
            in0 => \N__6773\,
            in1 => \N__8843\,
            in2 => \N__6812\,
            in3 => \N__6788\,
            lcout => \U712_CHIP_RAM.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__8795\,
            in2 => \N__8124\,
            in3 => \N__7841\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__8294\,
            in1 => \N__8796\,
            in2 => \N__8125\,
            in3 => \N__7241\,
            lcout => \U712_CHIP_RAM.CMA_5_3_ns_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101101011011"
        )
    port map (
            in0 => \N__8765\,
            in1 => \N__7757\,
            in2 => \N__8116\,
            in3 => \N__7829\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000001111"
        )
    port map (
            in0 => \N__7229\,
            in1 => \N__7214\,
            in2 => \N__7199\,
            in3 => \N__8766\,
            lcout => \U712_CHIP_RAM.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100111101"
        )
    port map (
            in0 => \N__7796\,
            in1 => \N__8764\,
            in2 => \N__8115\,
            in3 => \N__7835\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_5_3_ns_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000001111"
        )
    port map (
            in0 => \N__7187\,
            in1 => \N__7169\,
            in2 => \N__7148\,
            in3 => \N__8767\,
            lcout => \U712_CHIP_RAM.N_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__7751\,
            in1 => \N__7469\,
            in2 => \N__7134\,
            in3 => \N__7733\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9262\,
            ce => 'H',
            sr => \N__9037\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7078\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7628\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9267\,
            ce => 'H',
            sr => \N__9025\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7750\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9267\,
            ce => 'H',
            sr => \N__9025\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101000101"
        )
    port map (
            in0 => \N__7088\,
            in1 => \N__7592\,
            in2 => \N__7471\,
            in3 => \N__7074\,
            lcout => \CUMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011011111"
        )
    port map (
            in0 => \N__7461\,
            in1 => \N__7626\,
            in2 => \N__7596\,
            in3 => \N__7661\,
            lcout => \CLMBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111101"
        )
    port map (
            in0 => \N__7465\,
            in1 => \N__7627\,
            in2 => \N__7597\,
            in3 => \N__7544\,
            lcout => \CUUBEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.N_52_i_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7507\,
            in2 => \_gnd_net_\,
            in3 => \N__7472\,
            lcout => \N_52_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7384\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9240\,
            ce => \N__7956\,
            sr => \N__9076\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100011"
        )
    port map (
            in0 => \N__7346\,
            in1 => \N__8129\,
            in2 => \N__8473\,
            in3 => \N__8582\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9247\,
            ce => \N__8633\,
            sr => \N__9071\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_15_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__7319\,
            in1 => \_gnd_net_\,
            in2 => \N__8474\,
            in3 => \N__8581\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9247\,
            ce => \N__8633\,
            sr => \N__9071\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__7292\,
            in1 => \N__8342\,
            in2 => \N__9335\,
            in3 => \N__8839\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9247\,
            ce => \N__8633\,
            sr => \N__9071\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_8_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8180\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9256\,
            ce => \N__8266\,
            sr => \N__9063\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_6_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9256\,
            ce => \N__8266\,
            sr => \N__9063\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9263\,
            ce => \N__7941\,
            sr => \N__9056\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9263\,
            ce => \N__7941\,
            sr => \N__9056\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7823\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9263\,
            ce => \N__7941\,
            sr => \N__9056\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_1_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7816\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9268\,
            ce => \N__8250\,
            sr => \N__9044\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_2_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7790\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9268\,
            ce => \N__8250\,
            sr => \N__9044\
        );

    \U712_CHIP_RAM.CAS_SYNC_RNIB8S01_1_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__9118\,
            in1 => \N__7749\,
            in2 => \_gnd_net_\,
            in3 => \N__7732\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESS4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_0_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7717\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9277\,
            ce => \N__8251\,
            sr => \N__9026\
        );

    \U712_CHIP_RAM.RASn_LC_16_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8585\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9235\,
            ce => 'H',
            sr => \N__9080\
        );

    \U712_CHIP_RAM.WEn_LC_16_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8470\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9241\,
            ce => 'H',
            sr => \N__9079\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__8879\,
            in1 => \N__8341\,
            in2 => \N__8147\,
            in3 => \N__8840\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9250\,
            ce => \N__8654\,
            sr => \N__9077\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__8577\,
            in1 => \N__8117\,
            in2 => \_gnd_net_\,
            in3 => \N__8463\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_esr_4_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8323\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9264\,
            ce => \N__8279\,
            sr => \N__9068\
        );

    \CONSTANT_ONE_LUT4_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8176\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9269\,
            ce => \N__7931\,
            sr => \N__9072\
        );

    \U712_CHIP_RAM.CASn_LC_18_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8135\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9257\,
            ce => 'H',
            sr => \N__9081\
        );

    \U712_CHIP_RAM.RAS_SYNC_RNI9LBR_1_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__9121\,
            in1 => \N__7910\,
            in2 => \_gnd_net_\,
            in3 => \N__9298\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESS5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RAS_SYNC_1_LC_19_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9299\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9280\,
            ce => 'H',
            sr => \N__9078\
        );

    \U712_CHIP_RAM.RAS_SYNC_0_LC_19_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9328\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9308\,
            lcout => \U712_CHIP_RAM.RAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9280\,
            ce => 'H',
            sr => \N__9078\
        );
end \INTERFACE\;

----------------------------------------------------------------------------------
--This work is shared under the Attribution-NonCommercial-ShareAlike 4.0 International (CC BY-NC-SA 4.0) License
--https://creativecommons.org/licenses/by-nc-sa/4.0/legalcode
	
--You are free to:
--Share - copy and redistribute the material in any medium or format
--Adapt - remix, transform, and build upon the material

--Under the following terms:

--Attribution - You must give appropriate credit, provide a link to the license, and indicate if changes were made. 
--You may do so in any reasonable manner, but not in any way that suggests the licensor endorses you or your use.

--NonCommercial - You may not use the material for commercial purposes.

--ShareAlike - If you remix, transform, or build upon the material, you must distribute your contributions under the 
--same license as the original.

--No additional restrictions - You may not apply legal terms or technological measures that legally restrict others 
--from doing anything the license permits.
----------------------------------------------------------------------------------
-- Engineer:       JASON NEUS
-- 
-- Design Name:    AMIGA PCI U109
-- Project Name:   AMIGA PCI https://github.com/jasonsbeer/AmigaPCI
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PCI_CYCLE is

	Port ( 
	 
		A_HIGH : IN  STD_LOGIC_VECTOR (22 DOWNTO 20);
		A_LOW : IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		AD : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		BCLK : IN STD_LOGIC;
		PCICLK : IN STD_LOGIC;
		nRESET : IN STD_LOGIC;
		RnW : IN STD_LOGIC;
		nTS : IN STD_LOGIC;
		TT0 : IN STD_LOGIC;
		TT1 : IN STD_LOGIC;
		UPA0 : IN STD_LOGIC;
		UPA1 : IN STD_LOGIC;
		CPUSPACE : IN STD_LOGIC;
		BEN : IN STD_LOGIC;
		nDEVSEL : IN STD_LOGIC;
		nTRDY : IN STD_LOGIC;
		nSTOP : IN STD_LOGIC;
				
		nIRDY : INOUT STD_LOGIC;
		nFRAME : INOUT STD_LOGIC;
		CYCLE_DATA_PHASE : INOUT STD_LOGIC; --IDENTIFIES WHEN WE ARE IN A PCI CYCLE DATA PHASE.
		
		CPU_TRANSFER_ACK : OUT STD_LOGIC; --READY TO ASSERT _TA.
		CPU_TRANSFER_EACK : OUT STD_LOGIC; --READY TO ASSERT _TEA.
		PCI_TRANSFER_ACK_READY : OUT STD_LOGIC; --SETS PCI CYCLE TO ACTIVATE _TA SIGNAL.		
		AD_OUT : OUT STD_LOGIC_VECTOR (1 DOWNTO 0); --VECTOR TO MOVE AD BUS DATA FROM THE PROCESS TO THE PINS.
		nADDRESS_PHASE : OUT STD_LOGIC;
		AD_LATCH : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
		
			  
	);

end PCI_CYCLE;

architecture Behavioral of PCI_CYCLE is

	SIGNAL TRANSFER_START : STD_LOGIC; --LATCH THE START OF A NEW DATA TRANSFER CYCLE.
	SIGNAL TRANSFER_START_ACK : STD_LOGIC; --ACK THE START OF A NEW DATA TRANSFER CYCLE.
	SIGNAL BURST_CYCLE : STD_LOGIC; --ASSERT WHEN THE 68040 IS CALLING FOR A BURST TRANSFER.	
	SIGNAL CPU_TRANSFER_ACK_WAIT : STD_LOGIC_VECTOR (4 DOWNTO 0); --HOLD OFF ASSERTION OF _TA OR _TEA.
	SIGNAL PCI_TRANSFER_ACK : STD_LOGIC_VECTOR (3 DOWNTO 0); --HOLD OFF ASSERTION OF _TA OR _TEA.
	SIGNAL STOP_CYCLE : STD_LOGIC; --CONNECTED TO THE _STOP SIGNAL AND LATCHED ON THE RISING CLOCK EDGE.
	SIGNAL TARGET_READY : STD_LOGIC; --CONNECTED TO THE _TRDY SIGNAL AND LATCHED ON THE RISING CLOCK EDGE.
	SIGNAL DEVICE_SELECTED : STD_LOGIC; --THE TARGET DEVICE HAS ASSERTED _DEVSEL.	
	SIGNAL END_PCI_CYCLE : STD_LOGIC; --SIGNAL TO END THE PCI CYCLE AT THE END OF A BURST CYCLE
	SIGNAL RETRY_DISABLE : STD_LOGIC; --DISABLE RETRY CONDITIONS
	
	--THE TIMEOUT FOR A DEVICE TO ASSERT _DEVSEL.
	CONSTANT PCI_RESPONSE_TIMEOUT : INTEGER := 3; 
	SIGNAL PCI_RESPONSE_TIMEOUT_COUNT : INTEGER RANGE 0 TO PCI_RESPONSE_TIMEOUT;
	
	--TYPE PCI_STATE IS (IDLE, ADDRESS, DATA0, DATA1, DATA2, DATA3);
	TYPE PCI_STATE IS (IDLE, ADDRESS, DATA, TERMINATION);
	SIGNAL CURRENT_PCI_STATE : PCI_STATE;
	
	--THE NUMBER OF LONG WORDS IN A BURST CYCLE.
	CONSTANT PCI_BURST_COUNT : INTEGER := 3;
	SIGNAL PCI_DATA_PHASE : INTEGER RANGE 0 TO PCI_BURST_COUNT;
	
	--THE FOUR RECOGNIZED PCI BUS COMMANDS.
	TYPE PCI_AD_COMMAND IS (IO_SPACE, MEMORY_SPACE, CONFIG0_SPACE, CONFIG1_SPACE);
	SIGNAL CURRENT_PCI_COMMAND : PCI_AD_COMMAND;	

begin

	---------------------------------------
	-- MC68040 DATA TRANSFER START CYCLE --
	---------------------------------------

	--WE ASSERT THIS SIGNAL WHEN A NEW DATA TRANSFER CYCLE STARTS.
	--WHEN WE ACK THE START OF A NEW TRANSFER, THE SIGNAL IS RESET.
	--WE ALSO CAPTURE THE TRANSFER TYPE SIGNALS TO SEE IF THIS IS
	--A BURST TRANSFER AND DETERMINE THE APPROPRIATE PCI BUS COMMAND.
	--PROMETHEUS DRIVEN COMMANDS ARE QUALIFIED WITH THE BEN SIGNAL.
	
	BURST_CYCLE <= NOT TT0 AND TT1;

	PROCESS (BCLK, nRESET, TRANSFER_START_ACK) BEGIN
	
		IF nRESET = '0' OR TRANSFER_START_ACK = '1' THEN
		
			TRANSFER_START <= '0';
			--BURST_CYCLE <= '0';
			CURRENT_PCI_COMMAND <= MEMORY_SPACE;
		
		ELSIF RISING_EDGE (BCLK) THEN
		
			TRANSFER_START <= NOT CPUSPACE AND (NOT nTS OR TRANSFER_START);
			--BURST_CYCLE <= NOT TT0 AND TT1;
			
			IF BEN = '1' AND A_HIGH(22) = '1' AND A_HIGH(21) = '1' THEN
				CURRENT_PCI_COMMAND <= IO_SPACE;
			ELSIF (BEN = '1' AND A_HIGH(20) = '1') OR (UPA0 = '1' AND UPA1= '0') THEN
				CURRENT_PCI_COMMAND <= CONFIG1_SPACE;
			ELSIF (BEN = '1' AND A_HIGH(20) = '0') OR (UPA0 = '0' AND UPA1 = '0') THEN
				CURRENT_PCI_COMMAND <= CONFIG0_SPACE;
			ELSE
				CURRENT_PCI_COMMAND <= MEMORY_SPACE;
			END IF;
		
		END IF;	
	
	END PROCESS;		
	
	-------------------------------
	-- MC68040 DATA TRANSFER ACK --
	-------------------------------
	
	--CYCLE_DATA_PHASE <= '1' WHEN nGNT = '1' AND (CURRENT_PCI_STATE = DATA0 OR CURRENT_PCI_STATE = DATA1 OR CURRENT_PCI_STATE = DATA2 OR CURRENT_PCI_STATE = DATA3) ELSE '0';
	--CYCLE_DATA_PHASE <= '1' WHEN CURRENT_PCI_STATE = DATA0 OR CURRENT_PCI_STATE = DATA1 OR CURRENT_PCI_STATE = DATA2 OR CURRENT_PCI_STATE = DATA3 ELSE '0';
	CYCLE_DATA_PHASE <= '1' WHEN CURRENT_PCI_STATE = DATA ELSE '0';
	
	PCI_TRANSFER_ACK_READY <= CYCLE_DATA_PHASE OR NOT RETRY_DISABLE; -- RETRY_CONDITION; --PCI_RETRY_CYCLE;	
	--PCI_TRANSFER_ACK_READY <= '1' WHEN CURRENT_PCI_STATE = DATA OR PCI_RETRY_CYCLE = '1' ELSE '0';
	
	PROCESS (BCLK, nRESET) BEGIN
	
		IF nRESET = '0' THEN
		
			CPU_TRANSFER_ACK <= '0';
			CPU_TRANSFER_EACK <= '0';
			CPU_TRANSFER_ACK_WAIT <= (OTHERS => '0');
		
		ELSIF FALLING_EDGE(BCLK) THEN
		
			IF CURRENT_PCI_STATE = ADDRESS THEN
			
				CPU_TRANSFER_ACK_WAIT <= (OTHERS => '0');
				CPU_TRANSFER_EACK <= '0';
				CPU_TRANSFER_ACK <= '0';
		
			ELSIF CURRENT_PCI_STATE = TERMINATION THEN			
				
				IF CPU_TRANSFER_ACK_WAIT(4) = '0' THEN
					
					--ASSERT _TEA FOR ALL CONDITIONS.
					CPU_TRANSFER_EACK <= '1';
					CPU_TRANSFER_ACK_WAIT(4) <= '1';
					
					--ASSERT _TA FOR RETRY CONDITION ONLY.
					CPU_TRANSFER_ACK <= NOT RETRY_DISABLE; --RETRY_CONDITION;					
					
				ELSE
				
					CPU_TRANSFER_EACK <= '0';
					CPU_TRANSFER_ACK <= '0';
					
				END IF;
						
			ELSE		
				
				IF CPU_TRANSFER_ACK_WAIT(PCI_DATA_PHASE) = '0' AND PCI_TRANSFER_ACK(PCI_DATA_PHASE) = '1' THEN -- AND ((RnW = '1' AND TARGET_READY = '1') OR (RnW = '0' AND PCI_TRANSFER_ACK(PCI_DATA_PHASE) = '1')) THEN	
				
					CPU_TRANSFER_ACK <= '1';
					CPU_TRANSFER_ACK_WAIT(PCI_DATA_PHASE) <= '1'; --ONCE CPU_TRANSFER_ACK IS SET, WE CAN PROCEED WITH ASSERTING _IRDY.			
					
				ELSE
				
					CPU_TRANSFER_ACK <= '0';

				END IF;
			
			END IF;
		
		END IF;
	
	END PROCESS;	
	
	-----------------------------
	-- PCI CYCLE STATE MACHINE --
	-----------------------------
	
	--PCI SIGNALS ARE LATCHED ON THE RISING CLOCK EDGE, SO THIS IS WHERE MOST OF 
	--THE MEAT AND POTATOES ARE. DATA TRANSFER CONDITIONS ARE READ HERE TO MOVE
	--THE CYCLE FORWARD.
	
	PROCESS (PCICLK, nRESET) BEGIN
	
		IF nRESET = '0' THEN
		
			STOP_CYCLE <= '0';
			TARGET_READY <= '0';
			DEVICE_SELECTED <= '0';
			PCI_TRANSFER_ACK <= (OTHERS => '0');
			AD_LATCH <= (OTHERS => '0');
			PCI_RESPONSE_TIMEOUT_COUNT <= 0;
			RETRY_DISABLE  <= '0';
			PCI_DATA_PHASE <= 0;
			RETRY_DISABLE <= '0';
			
		ELSIF RISING_EDGE(PCICLK) THEN
		
			STOP_CYCLE <= NOT nSTOP; --SIGNAL LATCHED FOR PCI FALLING EDGE PROCESS
			TARGET_READY <= NOT nTRDY; --SIGNAL LATCHED FOR PCI FALLING EDGE PROCESS
			DEVICE_SELECTED <= NOT nDEVSEL; --SIGNAL LATCHED FOR PCI FALLING EDGE PROCESS
			RETRY_DISABLE <= (NOT RETRY_DISABLE AND NOT nTRDY) OR (RETRY_DISABLE AND NOT nDEVSEL); --DISABLES THE RETRY CONDITION AT THE FIRST ASSERTION OF _TRDY
			
			CASE CURRENT_PCI_STATE IS --STATE MACHINE STATES ARE SET IN THE FALLING EDGE PROCESS
			
				WHEN IDLE =>
			
					PCI_TRANSFER_ACK <= (OTHERS => '0'); --RESET VECTOR WHEN PCI STATE IS IDLE
					PCI_RESPONSE_TIMEOUT_COUNT <= 0; --RESET THE DEVICE RESPONSE TIMEOUT
					PCI_DATA_PHASE <= 0; --RESET THE BURST COUNTER
				
				WHEN ADDRESS =>
				
					IF nDEVSEL = '1' THEN PCI_RESPONSE_TIMEOUT_COUNT <= PCI_RESPONSE_TIMEOUT_COUNT + 1; END IF; --INCREMENT TIMEOUT COUNTER
					
				WHEN DATA =>
			
					IF nTRDY = '0' AND nSTOP = '1' THEN --AND PCI_TRANSFER_ACK(PCI_DATA_PHASE) = '0' THEN
					
						IF nIRDY = '0' THEN
							
							PCI_TRANSFER_ACK(PCI_DATA_PHASE) <= '1'; --SIGNAL PCI FALLING EDGE PROCESS TO NEGATE _IRDY
							IF RnW = '1' THEN AD_LATCH <= AD; END IF; --LATCH DATA FROM THE AD BUS ON READ CYCLES.
							
						ELSE
						
							PCI_DATA_PHASE <= PCI_DATA_PHASE + 1; --INCREMENT THE DATA PHASE BURST COUNTER
							
						END IF;
					
					END IF;		

				WHEN TERMINATION =>
				
			END CASE;
		
		END IF;
		
	END PROCESS;
	
	--WE DRIVE SIGNALS ON THE FALLING CLOCK EDGE HERE. THIS ENABLES COMMUNICATION WITH 
	--THE TARGET DEVICE BY ENSURING THE SIGNALS MEET SETUP TIMES FOR THE RISING EDGE SAMPLE.
	--DATA TRANSFER CONDITIONS ARE SET HERE TO MOVE THE CYCLE FORWARD.
	
	PROCESS (PCICLK, nRESET) BEGIN
	
		IF nRESET = '0' THEN
		
			CURRENT_PCI_STATE <= IDLE;
			TRANSFER_START_ACK <= '0';
			nFRAME <= '1';
			nADDRESS_PHASE <= '1';
			nIRDY <= '1';
			END_PCI_CYCLE <= '0';
		
		ELSIF FALLING_EDGE (PCICLK) THEN
		
			CASE CURRENT_PCI_STATE IS
			
				WHEN IDLE =>
				
					IF TRANSFER_START = '1' THEN --START THE PCI CYCLE!
						
						CURRENT_PCI_STATE <= ADDRESS;						
						TRANSFER_START_ACK <= '1';
						nFRAME <= '0';
						nADDRESS_PHASE <= '0';
						
						CASE CURRENT_PCI_COMMAND IS
						
							WHEN IO_SPACE =>
							
								AD_OUT <= A_LOW;
								--CBE <= "001" & NOT RnW;

							WHEN MEMORY_SPACE =>
							
								AD_OUT <= "1" & NOT BURST_CYCLE; --A(31 DOWNTO 2) & "1" & NOT BURST_CYCLE;
								--CBE <= "011" & NOT RnW;
							
							WHEN CONFIG0_SPACE =>
							
								AD_OUT <= "00"; --A(31 DOWNTO 2) & "00";
								--CBE <= "101" & NOT RnW;
							
							WHEN CONFIG1_SPACE =>
							
								AD_OUT <= "01"; --A(31 DOWNTO 2) & "01";
								--CBE <= "101" & NOT RnW;
							
						END CASE;							
					
					END IF;				
				
				WHEN ADDRESS =>
				
					nFRAME <= NOT BURST_CYCLE; --NEGATE _FRAME IF THIS IS NOT A BURST CYCLE
					TRANSFER_START_ACK <= '0'; --NEGATE TRANSFER START ACK
					nADDRESS_PHASE <= '1'; --NEGATE ADDRESS PHASE SIGNAL USED BY U110
					END_PCI_CYCLE <= '0'; --TURN OFF END PCI CYCLE SIGNAL
				
					IF DEVICE_SELECTED = '1' THEN
						
						IF STOP_CYCLE = '0' THEN
						
							CURRENT_PCI_STATE <= DATA;	
							nIRDY <= '0'; --ASSERT _IRDY BECAUSE WE ARE READY TO MOVE SOME DATA
							
						ELSE
						
							CURRENT_PCI_STATE <= TERMINATION;
							
						END IF;
							
					ELSE
					
						IF PCI_RESPONSE_TIMEOUT_COUNT = PCI_RESPONSE_TIMEOUT THEN
				
							nFRAME <= '1'; --NEGATE _FRAME ON BURST CYCLE BECAUSE NO DEVICE HAS REPLIED TO THE ADDRESS
							CURRENT_PCI_STATE <= IDLE;	----RETURN STATE MACHINE TO IDLE STATE BECUASE NO DEVICE CLAIMED THE CYCLE
						
						END IF;
					
					END IF;
				
				WHEN DATA =>
				
					IF STOP_CYCLE = '0' THEN
				
						nIRDY <= PCI_TRANSFER_ACK(PCI_DATA_PHASE); --SET _IRDY BASED ON WHERE WE ARE IN THIS DATA PHASE
					
						IF TARGET_READY = '1' THEN
						
							IF BURST_CYCLE = '1' THEN

								IF PCI_DATA_PHASE = PCI_BURST_COUNT THEN
									
									nFRAME <= '1'; --NEGATE FRAME BEFORE THE LAST DATA PHASE.
									END_PCI_CYCLE <= '1';								
								
								END IF;
								
								IF END_PCI_CYCLE = '1' THEN CURRENT_PCI_STATE <= IDLE; END IF; --RETURN STATE MACHINE TO IDLE STATE BECUASE TRANSFER IS DONE
								
							ELSE
							
								CURRENT_PCI_STATE <= IDLE; --RETURN STATE MACHINE TO IDLE STATE BECUASE TRANSFER IS DONE
							
							END IF;					
						
						END IF;
						
					ELSE
					
						CURRENT_PCI_STATE <= TERMINATION; --ACKNOWLEDGE THE END CYCLE REQUEST
						
					END IF;
				
				WHEN TERMINATION =>
				
					IF nIRDY = '1' THEN

						nFRAME <= '1'; --NEGATE FRAME BEFORE THE LAST DATA PHASE.
						nIRDY <= '0';
						
					ELSE
					
						nIRDY <= '1'; --NEGATE _IRDY
						CURRENT_PCI_STATE <= IDLE; --RETURN STATE MACHINE TO IDLE STATE BECUASE TRANSFER IS DONE
					
					END IF;
				
			END CASE;
		
		
		END IF;
		
	END PROCESS;
	

end Behavioral;
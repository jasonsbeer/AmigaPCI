-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 6 2025 19:31:10

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    TM : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : inout std_logic_vector(7 downto 4);
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    PIO_S0 : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    CIACS0n : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    PIO_P2 : out std_logic;
    CIACS1n : out std_logic;
    BRIDGE_ENn : out std_logic;
    PIO_S1 : out std_logic;
    ATA_MODE_S : in std_logic;
    PIO_P0 : out std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    REGSPACEn : out std_logic;
    TSn : in std_logic;
    RTC_ENn : out std_logic;
    PIO_S2 : out std_logic;
    ATA_ENn : out std_logic;
    TACKn : inout std_logic;
    ATA_MODE_P : in std_logic;
    ROMENn : out std_logic;
    PIO_P1 : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12497\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12404\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12386\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12368\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12341\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12332\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12323\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12305\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12287\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12260\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12251\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12224\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12179\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12142\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11824\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11442\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11257\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10950\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10944\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10890\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10768\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10730\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10568\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10345\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10280\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10229\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10223\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9440\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9417\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9276\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8737\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8241\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8127\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8019\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8010\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7973\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7863\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7848\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7839\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7659\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7344\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7266\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7236\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6930\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6549\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6387\ : std_logic;
signal \N__6384\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6234\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6065\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5799\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5685\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5112\ : std_logic;
signal \N__5109\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4998\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4728\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4384\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \PIO_S0_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \PIO_P0_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \U409_AUTOCONFIG.N_67_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_214_1\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_63\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_196_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_CONFC_net\ : std_logic;
signal \U409_AUTOCONFIG.ATA_BASE10Z0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.ATA_BASE10_cascade_\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_3\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_55_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.N_40\ : std_logic;
signal \U409_AUTOCONFIG.N_59_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_61\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_67\ : std_logic;
signal \U409_AUTOCONFIG.N_56\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0\ : std_logic;
signal \U409_AUTOCONFIG.N_59_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa\ : std_logic;
signal \U409_AUTOCONFIG.N_57\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\ : std_logic;
signal \AUTOCONFIG_SPACE_cascade_\ : std_logic;
signal \D_1_i\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_0\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_AZ0Z_18\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_a4Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTc_0_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_50\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTc_0_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_48\ : std_logic;
signal \U409_AUTOCONFIG.AC_START_RNI777KZ0Z2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG_D_OUT_0_i_2\ : std_logic;
signal \BRIDGE_BASE_1\ : std_logic;
signal \BRIDGE_BASE_2\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U409_AUTOCONFIG.N_68\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U409_AUTOCONFIG.N_47\ : std_logic;
signal \AUTOBOOT_c\ : std_logic;
signal \U409_AUTOCONFIG.N_196_1\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.N_54\ : std_logic;
signal \U409_ADDRESS_DECODE.g2_5_0\ : std_logic;
signal \U409_ADDRESS_DECODE.g2_6_0_cascade_\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_ADDRESS_DECODE.g2Z0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.g2Z0Z_10\ : std_logic;
signal \U409_ADDRESS_DECODE.g2Z0Z_11_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.g2Z0Z_9\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_1_0\ : std_logic;
signal \BRIDGE_BASE_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \ATA_BASE_5\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.g2Z0Z_5\ : std_logic;
signal \A_c_28\ : std_logic;
signal \U409_ADDRESS_DECODE_g2_6\ : std_logic;
signal \U409_ADDRESS_DECODE_g2_7_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_o7_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\ : std_logic;
signal \ATA_BASE_2\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_2C_net\ : std_logic;
signal \D_in_4\ : std_logic;
signal \D_in_5\ : std_logic;
signal \D_in_6\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\ : std_logic;
signal \BRIDGE_BASE_3\ : std_logic;
signal \un1_AUTOCONFIG_SPACE\ : std_logic;
signal \U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0\ : std_logic;
signal \D_in_7\ : std_logic;
signal \ATA_BASE_3\ : std_logic;
signal \INVU409_AUTOCONFIG.ATA_BASE_7C_net\ : std_logic;
signal \U409_ADDRESS_DECODE_ATA_ROM_d\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_0Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_o4Z0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE.g0_i_o4Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE_ATA_ROM_0_1\ : std_logic;
signal \U409_TRANSFER_ACK.CO1\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE.REG_SPACE_3\ : std_logic;
signal \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \A_c_17\ : std_logic;
signal \ATA_BASE_1\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_22\ : std_logic;
signal \ATA_BASE_0\ : std_logic;
signal \ATA_BASE_6\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_o7_2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_o7_4\ : std_logic;
signal \A_c_20\ : std_logic;
signal \ATA_BASE_7\ : std_logic;
signal \ATA_BASE_4\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_o7_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_13\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_TRANSFER_ACK.N_24\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_1_1\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_o7_6\ : std_logic;
signal \U409_TRANSFER_ACK.G_14_0_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.g0_0_0_o6_4\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\ : std_logic;
signal \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_ADDRESS_DECODE_ROMEN_1\ : std_logic;
signal \OVL_c\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \AUTOVECTOR\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_ADDRESS_DECODE_un2_REGSPACEn_0\ : std_logic;
signal \U409_ADDRESS_DECODE_Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_OUTnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_ATA_ROM_EN\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \U409_CIA.CLK_CIA6_4_cascade_\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_6_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\ : std_logic;
signal \bfn_12_9_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2\ : std_logic;
signal \U409_CIA.CLK_CIA6_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \bfn_14_5_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_14_8_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \PIO_P1_wire\ : std_logic;
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \ATA_MODE_P_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(1 downto 0);
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AUTOBOOT_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \PIO_P2_wire\ : std_logic;
signal \BRIDGE_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \PIO_P0_wire\ : std_logic;
signal \ATA_MODE_S_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \PIO_S0_wire\ : std_logic;
signal \PIO_S2_wire\ : std_logic;
signal \PIO_S1_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    PIO_P1 <= \PIO_P1_wire\;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \ATA_MODE_P_wire\ <= ATA_MODE_P;
    \TM_wire\ <= TM;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \AUTOBOOT_wire\ <= AUTOBOOT;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    PIO_P2 <= \PIO_P2_wire\;
    BRIDGE_ENn <= \BRIDGE_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    TICK60 <= \TICK60_wire\;
    PIO_P0 <= \PIO_P0_wire\;
    \ATA_MODE_S_wire\ <= ATA_MODE_S;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    BUFENn <= \BUFENn_wire\;
    PIO_S0 <= \PIO_S0_wire\;
    PIO_S2 <= \PIO_S2_wire\;
    PIO_S1 <= \PIO_S1_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__10297\,
            RESETB => \N__9759\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__12505\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12507\,
            DIN => \N__12506\,
            DOUT => \N__12505\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12507\,
            PADOUT => \N__12506\,
            PADIN => \N__12505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__12495\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12497\,
            DIN => \N__12496\,
            DOUT => \N__12495\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12497\,
            PADOUT => \N__12496\,
            PADIN => \N__12495\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__12485\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12487\,
            DIN => \N__12486\,
            DOUT => \N__12485\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12487\,
            PADOUT => \N__12486\,
            PADIN => \N__12485\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12476\,
            DIN => \N__12475\,
            DOUT => \N__12474\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12476\,
            PADOUT => \N__12475\,
            PADIN => \N__12474\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12467\,
            DIN => \N__12466\,
            DOUT => \N__12465\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12467\,
            PADOUT => \N__12466\,
            PADIN => \N__12465\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12458\,
            DIN => \N__12457\,
            DOUT => \N__12456\,
            PACKAGEPIN => \PIO_P1_wire\
        );

    \PIO_P1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12458\,
            PADOUT => \N__12457\,
            PADIN => \N__12456\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9786\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12449\,
            DIN => \N__12448\,
            DOUT => \N__12447\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12449\,
            PADOUT => \N__12448\,
            PADIN => \N__12447\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4861\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__4603\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12440\,
            DIN => \N__12439\,
            DOUT => \N__12438\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12440\,
            PADOUT => \N__12439\,
            PADIN => \N__12438\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12431\,
            DIN => \N__12430\,
            DOUT => \N__12429\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12431\,
            PADOUT => \N__12430\,
            PADIN => \N__12429\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12422\,
            DIN => \N__12421\,
            DOUT => \N__12420\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12422\,
            PADOUT => \N__12421\,
            PADIN => \N__12420\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6442\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12413\,
            DIN => \N__12412\,
            DOUT => \N__12411\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12413\,
            PADOUT => \N__12412\,
            PADIN => \N__12411\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_MODE_P_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12404\,
            DIN => \N__12403\,
            DOUT => \N__12402\,
            PACKAGEPIN => \ATA_MODE_P_wire\
        );

    \ATA_MODE_P_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12404\,
            PADOUT => \N__12403\,
            PADIN => \N__12402\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PIO_P0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12395\,
            DIN => \N__12394\,
            DOUT => \N__12393\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12395\,
            PADOUT => \N__12394\,
            PADIN => \N__12393\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4846\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__5020\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12386\,
            DIN => \N__12385\,
            DOUT => \N__12384\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12386\,
            PADOUT => \N__12385\,
            PADIN => \N__12384\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12377\,
            DIN => \N__12376\,
            DOUT => \N__12375\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12377\,
            PADOUT => \N__12376\,
            PADIN => \N__12375\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12368\,
            DIN => \N__12367\,
            DOUT => \N__12366\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12368\,
            PADOUT => \N__12367\,
            PADIN => \N__12366\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12359\,
            DIN => \N__12358\,
            DOUT => \N__12357\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12359\,
            PADOUT => \N__12358\,
            PADIN => \N__12357\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7681\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12350\,
            DIN => \N__12349\,
            DOUT => \N__12348\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12350\,
            PADOUT => \N__12349\,
            PADIN => \N__12348\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12341\,
            DIN => \N__12340\,
            DOUT => \N__12339\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12341\,
            PADOUT => \N__12340\,
            PADIN => \N__12339\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8833\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12332\,
            DIN => \N__12331\,
            DOUT => \N__12330\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12332\,
            PADOUT => \N__12331\,
            PADIN => \N__12330\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9874\,
            DIN0 => OPEN,
            DOUT0 => \N__9612\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AUTOBOOT_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12323\,
            DIN => \N__12322\,
            DOUT => \N__12321\,
            PACKAGEPIN => \AUTOBOOT_wire\
        );

    \AUTOBOOT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12323\,
            PADOUT => \N__12322\,
            PADIN => \N__12321\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AUTOBOOT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12314\,
            DIN => \N__12313\,
            DOUT => \N__12312\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12314\,
            PADOUT => \N__12313\,
            PADIN => \N__12312\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12305\,
            DIN => \N__12304\,
            DOUT => \N__12303\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12305\,
            PADOUT => \N__12304\,
            PADIN => \N__12303\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8290\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12296\,
            DIN => \N__12295\,
            DOUT => \N__12294\,
            PACKAGEPIN => \PIO_P2_wire\
        );

    \PIO_P2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12296\,
            PADOUT => \N__12295\,
            PADIN => \N__12294\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12287\,
            DIN => \N__12286\,
            DOUT => \N__12285\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12287\,
            PADOUT => \N__12286\,
            PADIN => \N__12285\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BRIDGE_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12278\,
            DIN => \N__12277\,
            DOUT => \N__12276\,
            PACKAGEPIN => \BRIDGE_ENn_wire\
        );

    \BRIDGE_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12278\,
            PADOUT => \N__12277\,
            PADIN => \N__12276\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6580\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12269\,
            DIN => \N__12268\,
            DOUT => \N__12267\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12269\,
            PADOUT => \N__12268\,
            PADIN => \N__12267\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12260\,
            DIN => \N__12259\,
            DOUT => \N__12258\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12260\,
            PADOUT => \N__12259\,
            PADIN => \N__12258\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12251\,
            DIN => \N__12250\,
            DOUT => \N__12249\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12251\,
            PADOUT => \N__12250\,
            PADIN => \N__12249\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12242\,
            DIN => \N__12241\,
            DOUT => \N__12240\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12242\,
            PADOUT => \N__12241\,
            PADIN => \N__12240\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12233\,
            DIN => \N__12232\,
            DOUT => \N__12231\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12233\,
            PADOUT => \N__12232\,
            PADIN => \N__12231\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9199\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12224\,
            DIN => \N__12223\,
            DOUT => \N__12222\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12224\,
            PADOUT => \N__12223\,
            PADIN => \N__12222\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10966\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12215\,
            DIN => \N__12214\,
            DOUT => \N__12213\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12215\,
            PADOUT => \N__12214\,
            PADIN => \N__12213\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12206\,
            DIN => \N__12205\,
            DOUT => \N__12204\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12206\,
            PADOUT => \N__12205\,
            PADIN => \N__12204\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4856\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__5050\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12197\,
            DIN => \N__12196\,
            DOUT => \N__12195\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12197\,
            PADOUT => \N__12196\,
            PADIN => \N__12195\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12188\,
            DIN => \N__12187\,
            DOUT => \N__12186\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12188\,
            PADOUT => \N__12187\,
            PADIN => \N__12186\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12179\,
            DIN => \N__12178\,
            DOUT => \N__12177\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12179\,
            PADOUT => \N__12178\,
            PADIN => \N__12177\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12170\,
            DIN => \N__12169\,
            DOUT => \N__12168\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12170\,
            PADOUT => \N__12169\,
            PADIN => \N__12168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6730\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12161\,
            DIN => \N__12160\,
            DOUT => \N__12159\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12161\,
            PADOUT => \N__12160\,
            PADIN => \N__12159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10621\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12152\,
            DIN => \N__12151\,
            DOUT => \N__12150\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12152\,
            PADOUT => \N__12151\,
            PADIN => \N__12150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_P0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12143\,
            DIN => \N__12142\,
            DOUT => \N__12141\,
            PACKAGEPIN => \PIO_P0_wire\
        );

    \PIO_P0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12143\,
            PADOUT => \N__12142\,
            PADIN => \N__12141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_MODE_S_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__12134\,
            DIN => \N__12133\,
            DOUT => \N__12132\,
            PACKAGEPIN => \ATA_MODE_S_wire\
        );

    \ATA_MODE_S_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12134\,
            PADOUT => \N__12133\,
            PADIN => \N__12132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PIO_S0_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12125\,
            DIN => \N__12124\,
            DOUT => \N__12123\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12125\,
            PADOUT => \N__12124\,
            PADIN => \N__12123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12116\,
            DIN => \N__12115\,
            DOUT => \N__12114\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12116\,
            PADOUT => \N__12115\,
            PADIN => \N__12114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9988\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12107\,
            DIN => \N__12106\,
            DOUT => \N__12105\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12107\,
            PADOUT => \N__12106\,
            PADIN => \N__12105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12098\,
            DIN => \N__12097\,
            DOUT => \N__12096\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12098\,
            PADOUT => \N__12097\,
            PADIN => \N__12096\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9154\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12089\,
            DIN => \N__12088\,
            DOUT => \N__12087\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12089\,
            PADOUT => \N__12088\,
            PADIN => \N__12087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12080\,
            DIN => \N__12079\,
            DOUT => \N__12078\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12080\,
            PADOUT => \N__12079\,
            PADIN => \N__12078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12071\,
            DIN => \N__12070\,
            DOUT => \N__12069\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12071\,
            PADOUT => \N__12070\,
            PADIN => \N__12069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10441\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12062\,
            DIN => \N__12061\,
            DOUT => \N__12060\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12062\,
            PADOUT => \N__12061\,
            PADIN => \N__12060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12053\,
            DIN => \N__12052\,
            DOUT => \N__12051\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12053\,
            PADOUT => \N__12052\,
            PADIN => \N__12051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9873\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__9600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12044\,
            DIN => \N__12043\,
            DOUT => \N__12042\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12044\,
            PADOUT => \N__12043\,
            PADIN => \N__12042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12035\,
            DIN => \N__12034\,
            DOUT => \N__12033\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12035\,
            PADOUT => \N__12034\,
            PADIN => \N__12033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9340\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12026\,
            DIN => \N__12025\,
            DOUT => \N__12024\,
            PACKAGEPIN => \PIO_S0_wire\
        );

    \PIO_S0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12026\,
            PADOUT => \N__12025\,
            PADIN => \N__12024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4444\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12017\,
            DIN => \N__12016\,
            DOUT => \N__12015\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12017\,
            PADOUT => \N__12016\,
            PADIN => \N__12015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12008\,
            DIN => \N__12007\,
            DOUT => \N__12006\,
            PACKAGEPIN => \PIO_S2_wire\
        );

    \PIO_S2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12008\,
            PADOUT => \N__12007\,
            PADIN => \N__12006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9799\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11999\,
            DIN => \N__11998\,
            DOUT => \N__11997\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11999\,
            PADOUT => \N__11998\,
            PADIN => \N__11997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4857\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__5872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11990\,
            DIN => \N__11989\,
            DOUT => \N__11988\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11990\,
            PADOUT => \N__11989\,
            PADIN => \N__11988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11981\,
            DIN => \N__11980\,
            DOUT => \N__11979\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11981\,
            PADOUT => \N__11980\,
            PADIN => \N__11979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PIO_S1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11972\,
            DIN => \N__11971\,
            DOUT => \N__11970\,
            PACKAGEPIN => \PIO_S1_wire\
        );

    \PIO_S1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11972\,
            PADOUT => \N__11971\,
            PADIN => \N__11970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11963\,
            DIN => \N__11962\,
            DOUT => \N__11961\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11963\,
            PADOUT => \N__11962\,
            PADIN => \N__11961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11954\,
            DIN => \N__11953\,
            DOUT => \N__11952\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11954\,
            PADOUT => \N__11953\,
            PADIN => \N__11952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11945\,
            DIN => \N__11944\,
            DOUT => \N__11943\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11945\,
            PADOUT => \N__11944\,
            PADIN => \N__11943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11936\,
            DIN => \N__11935\,
            DOUT => \N__11934\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11936\,
            PADOUT => \N__11935\,
            PADIN => \N__11934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11927\,
            DIN => \N__11926\,
            DOUT => \N__11925\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11927\,
            PADOUT => \N__11926\,
            PADIN => \N__11925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11918\,
            DIN => \N__11917\,
            DOUT => \N__11916\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11918\,
            PADOUT => \N__11917\,
            PADIN => \N__11916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11909\,
            DIN => \N__11908\,
            DOUT => \N__11907\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11909\,
            PADOUT => \N__11908\,
            PADIN => \N__11907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9823\,
            DIN0 => OPEN,
            DOUT0 => \N__9613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2885\ : InMux
    port map (
            O => \N__11890\,
            I => \N__11886\
        );

    \I__2884\ : InMux
    port map (
            O => \N__11889\,
            I => \N__11883\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__11886\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2882\ : LocalMux
    port map (
            O => \N__11883\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2881\ : InMux
    port map (
            O => \N__11878\,
            I => \N__11875\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__11875\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2879\ : InMux
    port map (
            O => \N__11872\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2878\ : InMux
    port map (
            O => \N__11869\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2877\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11862\
        );

    \I__2876\ : InMux
    port map (
            O => \N__11865\,
            I => \N__11859\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__11862\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__11859\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2873\ : ClkMux
    port map (
            O => \N__11854\,
            I => \N__11827\
        );

    \I__2872\ : ClkMux
    port map (
            O => \N__11853\,
            I => \N__11827\
        );

    \I__2871\ : ClkMux
    port map (
            O => \N__11852\,
            I => \N__11827\
        );

    \I__2870\ : ClkMux
    port map (
            O => \N__11851\,
            I => \N__11827\
        );

    \I__2869\ : ClkMux
    port map (
            O => \N__11850\,
            I => \N__11827\
        );

    \I__2868\ : ClkMux
    port map (
            O => \N__11849\,
            I => \N__11827\
        );

    \I__2867\ : ClkMux
    port map (
            O => \N__11848\,
            I => \N__11827\
        );

    \I__2866\ : ClkMux
    port map (
            O => \N__11847\,
            I => \N__11827\
        );

    \I__2865\ : ClkMux
    port map (
            O => \N__11846\,
            I => \N__11827\
        );

    \I__2864\ : GlobalMux
    port map (
            O => \N__11827\,
            I => \N__11824\
        );

    \I__2863\ : gio2CtrlBuf
    port map (
            O => \N__11824\,
            I => \CLK6_c_g\
        );

    \I__2862\ : InMux
    port map (
            O => \N__11821\,
            I => \N__11817\
        );

    \I__2861\ : InMux
    port map (
            O => \N__11820\,
            I => \N__11814\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__11817\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2859\ : LocalMux
    port map (
            O => \N__11814\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2858\ : InMux
    port map (
            O => \N__11809\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2857\ : InMux
    port map (
            O => \N__11806\,
            I => \N__11802\
        );

    \I__2856\ : InMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__2855\ : LocalMux
    port map (
            O => \N__11802\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__11799\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2853\ : InMux
    port map (
            O => \N__11794\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2852\ : InMux
    port map (
            O => \N__11791\,
            I => \N__11787\
        );

    \I__2851\ : InMux
    port map (
            O => \N__11790\,
            I => \N__11784\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__11787\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__11784\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11779\,
            I => \N__11776\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__11776\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2846\ : InMux
    port map (
            O => \N__11773\,
            I => \bfn_14_8_0_\
        );

    \I__2845\ : InMux
    port map (
            O => \N__11770\,
            I => \N__11766\
        );

    \I__2844\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__11766\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__11763\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2841\ : InMux
    port map (
            O => \N__11758\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__11755\,
            I => \N__11752\
        );

    \I__2839\ : InMux
    port map (
            O => \N__11752\,
            I => \N__11748\
        );

    \I__2838\ : InMux
    port map (
            O => \N__11751\,
            I => \N__11745\
        );

    \I__2837\ : LocalMux
    port map (
            O => \N__11748\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11745\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2835\ : InMux
    port map (
            O => \N__11740\,
            I => \N__11737\
        );

    \I__2834\ : LocalMux
    port map (
            O => \N__11737\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2833\ : InMux
    port map (
            O => \N__11734\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2832\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11727\
        );

    \I__2831\ : InMux
    port map (
            O => \N__11730\,
            I => \N__11724\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11727\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__11724\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2828\ : InMux
    port map (
            O => \N__11719\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2827\ : InMux
    port map (
            O => \N__11716\,
            I => \N__11712\
        );

    \I__2826\ : InMux
    port map (
            O => \N__11715\,
            I => \N__11709\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__11712\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2824\ : LocalMux
    port map (
            O => \N__11709\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2823\ : InMux
    port map (
            O => \N__11704\,
            I => \N__11701\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__11701\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2821\ : InMux
    port map (
            O => \N__11698\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11691\
        );

    \I__2819\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__11691\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__11688\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11683\,
            I => \N__11680\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__11680\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11677\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2813\ : InMux
    port map (
            O => \N__11674\,
            I => \N__11670\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11673\,
            I => \N__11667\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__11670\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2810\ : LocalMux
    port map (
            O => \N__11667\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2809\ : InMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11659\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2807\ : InMux
    port map (
            O => \N__11656\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__2806\ : InMux
    port map (
            O => \N__11653\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__2805\ : InMux
    port map (
            O => \N__11650\,
            I => \N__11646\
        );

    \I__2804\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11643\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__11646\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__11643\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \N__11634\
        );

    \I__2800\ : InMux
    port map (
            O => \N__11637\,
            I => \N__11628\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11634\,
            I => \N__11628\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11633\,
            I => \N__11625\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__11628\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__11625\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__2794\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11611\
        );

    \I__2793\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11606\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11606\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11614\,
            I => \N__11603\
        );

    \I__2790\ : LocalMux
    port map (
            O => \N__11611\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11606\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__11603\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2787\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11592\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11595\,
            I => \N__11589\
        );

    \I__2785\ : LocalMux
    port map (
            O => \N__11592\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__11589\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11584\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2782\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11577\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11580\,
            I => \N__11574\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__11577\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2779\ : LocalMux
    port map (
            O => \N__11574\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2778\ : InMux
    port map (
            O => \N__11569\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2777\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11562\
        );

    \I__2776\ : InMux
    port map (
            O => \N__11565\,
            I => \N__11559\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__11562\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11559\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2773\ : InMux
    port map (
            O => \N__11554\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__2771\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11544\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11547\,
            I => \N__11541\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11544\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11541\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2767\ : CascadeMux
    port map (
            O => \N__11536\,
            I => \N__11533\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11530\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11527\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2763\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__2762\ : LocalMux
    port map (
            O => \N__11521\,
            I => \N__11517\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11520\,
            I => \N__11514\
        );

    \I__2760\ : Odrv4
    port map (
            O => \N__11517\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__11514\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__2757\ : InMux
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11503\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2755\ : InMux
    port map (
            O => \N__11500\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2754\ : InMux
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__11494\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11491\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__2751\ : InMux
    port map (
            O => \N__11488\,
            I => \N__11484\
        );

    \I__2750\ : InMux
    port map (
            O => \N__11487\,
            I => \N__11481\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__11484\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__11481\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2747\ : InMux
    port map (
            O => \N__11476\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11473\,
            I => \N__11469\
        );

    \I__2745\ : InMux
    port map (
            O => \N__11472\,
            I => \N__11466\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__11469\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__11466\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__2741\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11455\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__11455\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11452\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__2738\ : InMux
    port map (
            O => \N__11449\,
            I => \N__11445\
        );

    \I__2737\ : InMux
    port map (
            O => \N__11448\,
            I => \N__11442\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__11445\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11442\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__2733\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11431\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__11431\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2731\ : InMux
    port map (
            O => \N__11428\,
            I => \bfn_14_6_0_\
        );

    \I__2730\ : InMux
    port map (
            O => \N__11425\,
            I => \N__11421\
        );

    \I__2729\ : InMux
    port map (
            O => \N__11424\,
            I => \N__11418\
        );

    \I__2728\ : LocalMux
    port map (
            O => \N__11421\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__11418\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2726\ : InMux
    port map (
            O => \N__11413\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__2725\ : InMux
    port map (
            O => \N__11410\,
            I => \N__11406\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11409\,
            I => \N__11403\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__11406\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__11403\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2721\ : InMux
    port map (
            O => \N__11398\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__2720\ : InMux
    port map (
            O => \N__11395\,
            I => \N__11391\
        );

    \I__2719\ : InMux
    port map (
            O => \N__11394\,
            I => \N__11388\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__11391\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__11388\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11383\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11376\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11373\
        );

    \I__2713\ : LocalMux
    port map (
            O => \N__11376\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2712\ : LocalMux
    port map (
            O => \N__11373\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2711\ : InMux
    port map (
            O => \N__11368\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__2710\ : CascadeMux
    port map (
            O => \N__11365\,
            I => \N__11362\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11362\,
            I => \N__11358\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11361\,
            I => \N__11355\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11358\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11355\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11350\,
            I => \N__11347\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__11347\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2703\ : InMux
    port map (
            O => \N__11344\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__2702\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11338\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11338\,
            I => \U409_TICK.TICK503_11\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__11335\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__11332\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__11329\,
            I => \N__11325\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11328\,
            I => \N__11316\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11325\,
            I => \N__11307\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11324\,
            I => \N__11307\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11323\,
            I => \N__11307\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11322\,
            I => \N__11307\
        );

    \I__2692\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11300\
        );

    \I__2691\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11300\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11300\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11316\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__11307\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2687\ : LocalMux
    port map (
            O => \N__11300\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2686\ : InMux
    port map (
            O => \N__11293\,
            I => \N__11283\
        );

    \I__2685\ : InMux
    port map (
            O => \N__11292\,
            I => \N__11274\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11274\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11290\,
            I => \N__11274\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11289\,
            I => \N__11274\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11288\,
            I => \N__11267\
        );

    \I__2680\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11267\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11286\,
            I => \N__11267\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11283\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11274\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__11267\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__11260\,
            I => \N__11254\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__11259\,
            I => \N__11250\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__11258\,
            I => \N__11244\
        );

    \I__2672\ : InMux
    port map (
            O => \N__11257\,
            I => \N__11241\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11254\,
            I => \N__11236\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11253\,
            I => \N__11236\
        );

    \I__2669\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11233\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11249\,
            I => \N__11224\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11248\,
            I => \N__11224\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11224\
        );

    \I__2665\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11224\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11241\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__11236\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11233\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11224\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11215\,
            I => \N__11211\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11214\,
            I => \N__11207\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11211\,
            I => \N__11204\
        );

    \I__2657\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11201\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11207\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2655\ : Odrv4
    port map (
            O => \N__11204\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__11201\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2653\ : CascadeMux
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11185\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11180\
        );

    \I__2650\ : InMux
    port map (
            O => \N__11191\,
            I => \N__11180\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11188\,
            I => \N__11177\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__11185\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11180\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11177\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2645\ : CascadeMux
    port map (
            O => \N__11170\,
            I => \N__11167\
        );

    \I__2644\ : InMux
    port map (
            O => \N__11167\,
            I => \N__11163\
        );

    \I__2643\ : InMux
    port map (
            O => \N__11166\,
            I => \N__11160\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__11163\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11160\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2640\ : InMux
    port map (
            O => \N__11155\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__2639\ : InMux
    port map (
            O => \N__11152\,
            I => \N__11148\
        );

    \I__2638\ : InMux
    port map (
            O => \N__11151\,
            I => \N__11145\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__11148\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__11145\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2635\ : InMux
    port map (
            O => \N__11140\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__2634\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11133\
        );

    \I__2633\ : InMux
    port map (
            O => \N__11136\,
            I => \N__11130\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__11133\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__11130\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11125\,
            I => \N__11122\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__11122\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2628\ : InMux
    port map (
            O => \N__11119\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__2627\ : CascadeMux
    port map (
            O => \N__11116\,
            I => \N__11113\
        );

    \I__2626\ : InMux
    port map (
            O => \N__11113\,
            I => \N__11109\
        );

    \I__2625\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11106\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__11109\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__11106\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2622\ : InMux
    port map (
            O => \N__11101\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__2621\ : InMux
    port map (
            O => \N__11098\,
            I => \N__11094\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11097\,
            I => \N__11091\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__11094\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11091\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__11086\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__11083\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__11077\,
            I => \N__11070\
        );

    \I__2613\ : InMux
    port map (
            O => \N__11076\,
            I => \N__11059\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11059\
        );

    \I__2611\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11059\
        );

    \I__2610\ : InMux
    port map (
            O => \N__11073\,
            I => \N__11059\
        );

    \I__2609\ : InMux
    port map (
            O => \N__11070\,
            I => \N__11052\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11069\,
            I => \N__11052\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11052\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__11059\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11052\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2604\ : CascadeMux
    port map (
            O => \N__11047\,
            I => \N__11038\
        );

    \I__2603\ : CascadeMux
    port map (
            O => \N__11046\,
            I => \N__11035\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11045\,
            I => \N__11032\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11044\,
            I => \N__11025\
        );

    \I__2600\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11025\
        );

    \I__2599\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11025\
        );

    \I__2598\ : InMux
    port map (
            O => \N__11041\,
            I => \N__11018\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11038\,
            I => \N__11018\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11035\,
            I => \N__11018\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11032\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11025\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__11018\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2592\ : CascadeMux
    port map (
            O => \N__11011\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__2591\ : InMux
    port map (
            O => \N__11008\,
            I => \N__11005\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__11005\,
            I => \U409_TICK.TICK603_11\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__11002\,
            I => \N__10999\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10999\,
            I => \N__10989\
        );

    \I__2587\ : InMux
    port map (
            O => \N__10998\,
            I => \N__10982\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10997\,
            I => \N__10982\
        );

    \I__2585\ : InMux
    port map (
            O => \N__10996\,
            I => \N__10982\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10973\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10973\
        );

    \I__2582\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10973\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10973\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__10989\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__10982\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10973\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2577\ : IoInMux
    port map (
            O => \N__10966\,
            I => \N__10963\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10963\,
            I => \N__10960\
        );

    \I__2575\ : Span12Mux_s0_v
    port map (
            O => \N__10960\,
            I => \N__10957\
        );

    \I__2574\ : Span12Mux_v
    port map (
            O => \N__10957\,
            I => \N__10953\
        );

    \I__2573\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10950\
        );

    \I__2572\ : Odrv12
    port map (
            O => \N__10953\,
            I => \TICK50_c\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10950\,
            I => \TICK50_c\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10945\,
            I => \N__10937\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10944\,
            I => \N__10937\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10943\,
            I => \N__10932\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10932\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10937\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10932\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10919\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10926\,
            I => \N__10919\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10925\,
            I => \N__10914\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10914\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10919\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__10914\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__10909\,
            I => \N__10904\
        );

    \I__2557\ : CascadeMux
    port map (
            O => \N__10908\,
            I => \N__10900\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10907\,
            I => \N__10895\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10895\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10890\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10900\,
            I => \N__10890\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10895\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10890\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__10885\,
            I => \N__10877\
        );

    \I__2549\ : InMux
    port map (
            O => \N__10884\,
            I => \N__10874\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10883\,
            I => \N__10871\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10882\,
            I => \N__10866\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10866\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10880\,
            I => \N__10861\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10861\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__10874\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__10871\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10866\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__10861\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10848\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10845\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10848\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10845\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__2535\ : InMux
    port map (
            O => \N__10840\,
            I => \N__10837\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10837\,
            I => \N__10829\
        );

    \I__2533\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10826\
        );

    \I__2532\ : CascadeMux
    port map (
            O => \N__10835\,
            I => \N__10819\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__10834\,
            I => \N__10816\
        );

    \I__2530\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10813\
        );

    \I__2529\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10810\
        );

    \I__2528\ : Span4Mux_v
    port map (
            O => \N__10829\,
            I => \N__10803\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__10826\,
            I => \N__10803\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10825\,
            I => \N__10796\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10824\,
            I => \N__10796\
        );

    \I__2524\ : InMux
    port map (
            O => \N__10823\,
            I => \N__10796\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10822\,
            I => \N__10793\
        );

    \I__2522\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10788\
        );

    \I__2521\ : InMux
    port map (
            O => \N__10816\,
            I => \N__10788\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10783\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10783\
        );

    \I__2518\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10780\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__10808\,
            I => \N__10777\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__10803\,
            I => \N__10773\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10768\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__10793\,
            I => \N__10768\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__10788\,
            I => \N__10764\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__10783\,
            I => \N__10759\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__10780\,
            I => \N__10759\
        );

    \I__2510\ : InMux
    port map (
            O => \N__10777\,
            I => \N__10756\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10776\,
            I => \N__10753\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__10773\,
            I => \N__10746\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__10768\,
            I => \N__10746\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10767\,
            I => \N__10742\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__10764\,
            I => \N__10730\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__10759\,
            I => \N__10730\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10730\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10753\,
            I => \N__10730\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10752\,
            I => \N__10725\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10751\,
            I => \N__10725\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__10746\,
            I => \N__10721\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10718\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__10742\,
            I => \N__10715\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10741\,
            I => \N__10711\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10708\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10739\,
            I => \N__10705\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10730\,
            I => \N__10702\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10725\,
            I => \N__10699\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10696\
        );

    \I__2490\ : Span4Mux_h
    port map (
            O => \N__10721\,
            I => \N__10692\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10718\,
            I => \N__10689\
        );

    \I__2488\ : Span4Mux_h
    port map (
            O => \N__10715\,
            I => \N__10686\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10714\,
            I => \N__10683\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10676\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10676\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__10705\,
            I => \N__10676\
        );

    \I__2483\ : Span4Mux_h
    port map (
            O => \N__10702\,
            I => \N__10669\
        );

    \I__2482\ : Span4Mux_h
    port map (
            O => \N__10699\,
            I => \N__10669\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10696\,
            I => \N__10669\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10695\,
            I => \N__10666\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__10692\,
            I => \N__10663\
        );

    \I__2478\ : Span12Mux_s11_v
    port map (
            O => \N__10689\,
            I => \N__10656\
        );

    \I__2477\ : Sp12to4
    port map (
            O => \N__10686\,
            I => \N__10656\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10683\,
            I => \N__10656\
        );

    \I__2475\ : Span4Mux_v
    port map (
            O => \N__10676\,
            I => \N__10649\
        );

    \I__2474\ : Span4Mux_v
    port map (
            O => \N__10669\,
            I => \N__10649\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10649\
        );

    \I__2472\ : Sp12to4
    port map (
            O => \N__10663\,
            I => \N__10642\
        );

    \I__2471\ : Span12Mux_v
    port map (
            O => \N__10656\,
            I => \N__10642\
        );

    \I__2470\ : Sp12to4
    port map (
            O => \N__10649\,
            I => \N__10642\
        );

    \I__2469\ : Span12Mux_h
    port map (
            O => \N__10642\,
            I => \N__10639\
        );

    \I__2468\ : Odrv12
    port map (
            O => \N__10639\,
            I => \RESETn_c\
        );

    \I__2467\ : IoInMux
    port map (
            O => \N__10636\,
            I => \N__10633\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10630\
        );

    \I__2465\ : Span12Mux_s2_v
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__2464\ : Odrv12
    port map (
            O => \N__10627\,
            I => \RESETn_c_i\
        );

    \I__2463\ : CascadeMux
    port map (
            O => \N__10624\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__2462\ : IoInMux
    port map (
            O => \N__10621\,
            I => \N__10618\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__10618\,
            I => \N__10615\
        );

    \I__2460\ : Span4Mux_s3_v
    port map (
            O => \N__10615\,
            I => \N__10612\
        );

    \I__2459\ : Span4Mux_v
    port map (
            O => \N__10612\,
            I => \N__10609\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__10609\,
            I => \N__10605\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10602\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__10605\,
            I => \TICK60_c\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__10602\,
            I => \TICK60_c\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10597\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10594\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10588\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10588\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10585\,
            I => \N__10582\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10582\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10579\,
            I => \N__10574\
        );

    \I__2447\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10571\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10577\,
            I => \N__10568\
        );

    \I__2445\ : LocalMux
    port map (
            O => \N__10574\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10571\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__10568\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__2442\ : CascadeMux
    port map (
            O => \N__10561\,
            I => \N__10557\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10553\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10550\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10547\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10553\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10550\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10547\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__10540\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10529\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10536\,
            I => \N__10524\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10524\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10519\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10519\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10532\,
            I => \N__10516\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__10529\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10524\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10519\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10516\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10507\,
            I => \N__10504\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__10504\,
            I => \U409_CIA.CIA_CLK_COUNT11_2\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__2420\ : InMux
    port map (
            O => \N__10497\,
            I => \N__10492\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10492\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__10489\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_cascade_\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10486\,
            I => \N__10483\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__10483\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\
        );

    \I__2415\ : ClkMux
    port map (
            O => \N__10480\,
            I => \N__10468\
        );

    \I__2414\ : ClkMux
    port map (
            O => \N__10479\,
            I => \N__10468\
        );

    \I__2413\ : ClkMux
    port map (
            O => \N__10478\,
            I => \N__10468\
        );

    \I__2412\ : ClkMux
    port map (
            O => \N__10477\,
            I => \N__10468\
        );

    \I__2411\ : GlobalMux
    port map (
            O => \N__10468\,
            I => \N__10465\
        );

    \I__2410\ : gio2CtrlBuf
    port map (
            O => \N__10465\,
            I => \CLK28_IN_c_g\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10462\,
            I => \N__10456\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10451\
        );

    \I__2407\ : InMux
    port map (
            O => \N__10460\,
            I => \N__10451\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10448\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10456\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10451\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10448\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__2402\ : IoInMux
    port map (
            O => \N__10441\,
            I => \N__10438\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10438\,
            I => \N__10435\
        );

    \I__2400\ : Span4Mux_s2_v
    port map (
            O => \N__10435\,
            I => \N__10432\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__10432\,
            I => \N__10428\
        );

    \I__2398\ : InMux
    port map (
            O => \N__10431\,
            I => \N__10425\
        );

    \I__2397\ : Span4Mux_v
    port map (
            O => \N__10428\,
            I => \N__10421\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10425\,
            I => \N__10418\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10414\
        );

    \I__2394\ : Sp12to4
    port map (
            O => \N__10421\,
            I => \N__10409\
        );

    \I__2393\ : Span12Mux_h
    port map (
            O => \N__10418\,
            I => \N__10409\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10404\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10404\
        );

    \I__2390\ : Odrv12
    port map (
            O => \N__10409\,
            I => \CLK_CIA_c\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__10404\,
            I => \CLK_CIA_c\
        );

    \I__2388\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10396\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10396\,
            I => \U409_CIA.CLK_CIA_r_1_0\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__10393\,
            I => \N__10384\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10392\,
            I => \N__10381\
        );

    \I__2384\ : InMux
    port map (
            O => \N__10391\,
            I => \N__10376\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10390\,
            I => \N__10376\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10389\,
            I => \N__10373\
        );

    \I__2381\ : InMux
    port map (
            O => \N__10388\,
            I => \N__10370\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10387\,
            I => \N__10367\
        );

    \I__2379\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10364\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10381\,
            I => \N__10360\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__10376\,
            I => \N__10353\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10373\,
            I => \N__10345\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10370\,
            I => \N__10342\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10339\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10364\,
            I => \N__10336\
        );

    \I__2372\ : ClkMux
    port map (
            O => \N__10363\,
            I => \N__10303\
        );

    \I__2371\ : Glb2LocalMux
    port map (
            O => \N__10360\,
            I => \N__10303\
        );

    \I__2370\ : ClkMux
    port map (
            O => \N__10359\,
            I => \N__10303\
        );

    \I__2369\ : ClkMux
    port map (
            O => \N__10358\,
            I => \N__10303\
        );

    \I__2368\ : ClkMux
    port map (
            O => \N__10357\,
            I => \N__10303\
        );

    \I__2367\ : ClkMux
    port map (
            O => \N__10356\,
            I => \N__10303\
        );

    \I__2366\ : Glb2LocalMux
    port map (
            O => \N__10353\,
            I => \N__10303\
        );

    \I__2365\ : ClkMux
    port map (
            O => \N__10352\,
            I => \N__10303\
        );

    \I__2364\ : ClkMux
    port map (
            O => \N__10351\,
            I => \N__10303\
        );

    \I__2363\ : ClkMux
    port map (
            O => \N__10350\,
            I => \N__10303\
        );

    \I__2362\ : ClkMux
    port map (
            O => \N__10349\,
            I => \N__10303\
        );

    \I__2361\ : ClkMux
    port map (
            O => \N__10348\,
            I => \N__10303\
        );

    \I__2360\ : Glb2LocalMux
    port map (
            O => \N__10345\,
            I => \N__10303\
        );

    \I__2359\ : Glb2LocalMux
    port map (
            O => \N__10342\,
            I => \N__10303\
        );

    \I__2358\ : Glb2LocalMux
    port map (
            O => \N__10339\,
            I => \N__10303\
        );

    \I__2357\ : Glb2LocalMux
    port map (
            O => \N__10336\,
            I => \N__10303\
        );

    \I__2356\ : GlobalMux
    port map (
            O => \N__10303\,
            I => \N__10300\
        );

    \I__2355\ : gio2CtrlBuf
    port map (
            O => \N__10300\,
            I => \CLK40_IN_c_g\
        );

    \I__2354\ : IoInMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__10294\,
            I => \N__10291\
        );

    \I__2352\ : Span12Mux_s6_v
    port map (
            O => \N__10291\,
            I => \N__10288\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__10288\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10285\,
            I => \N__10280\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10284\,
            I => \N__10275\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10283\,
            I => \N__10275\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10280\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10275\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10264\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10261\
        );

    \I__2343\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10256\
        );

    \I__2342\ : InMux
    port map (
            O => \N__10267\,
            I => \N__10256\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10264\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10261\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__10256\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10249\,
            I => \N__10245\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10248\,
            I => \N__10242\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__10245\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10242\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__2334\ : CascadeMux
    port map (
            O => \N__10237\,
            I => \N__10234\
        );

    \I__2333\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10231\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10226\
        );

    \I__2331\ : InMux
    port map (
            O => \N__10230\,
            I => \N__10223\
        );

    \I__2330\ : InMux
    port map (
            O => \N__10229\,
            I => \N__10220\
        );

    \I__2329\ : Span4Mux_v
    port map (
            O => \N__10226\,
            I => \N__10217\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__10223\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10220\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__10217\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__10210\,
            I => \U409_TRANSFER_ACK.N_6_0_cascade_\
        );

    \I__2324\ : InMux
    port map (
            O => \N__10207\,
            I => \N__10204\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__10203\,
            I => \N__10195\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__10202\,
            I => \N__10192\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__10201\,
            I => \N__10188\
        );

    \I__2319\ : Span4Mux_h
    port map (
            O => \N__10198\,
            I => \N__10185\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10195\,
            I => \N__10180\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10180\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10191\,
            I => \N__10175\
        );

    \I__2315\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10175\
        );

    \I__2314\ : Odrv4
    port map (
            O => \N__10185\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10180\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10175\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2311\ : InMux
    port map (
            O => \N__10168\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10165\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10162\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10159\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__2307\ : CascadeMux
    port map (
            O => \N__10156\,
            I => \N__10152\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10149\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10152\,
            I => \N__10146\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__10149\,
            I => \N__10143\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10146\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__10143\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__10138\,
            I => \N__10135\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10126\
        );

    \I__2299\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10126\
        );

    \I__2298\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10123\
        );

    \I__2297\ : InMux
    port map (
            O => \N__10132\,
            I => \N__10118\
        );

    \I__2296\ : InMux
    port map (
            O => \N__10131\,
            I => \N__10118\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__10126\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10123\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10118\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__2292\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10107\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10101\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10107\,
            I => \N__10098\
        );

    \I__2289\ : InMux
    port map (
            O => \N__10106\,
            I => \N__10093\
        );

    \I__2288\ : InMux
    port map (
            O => \N__10105\,
            I => \N__10093\
        );

    \I__2287\ : InMux
    port map (
            O => \N__10104\,
            I => \N__10090\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__10101\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__10098\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10093\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10090\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__2282\ : SRMux
    port map (
            O => \N__10081\,
            I => \N__10077\
        );

    \I__2281\ : SRMux
    port map (
            O => \N__10080\,
            I => \N__10073\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10077\,
            I => \N__10070\
        );

    \I__2279\ : SRMux
    port map (
            O => \N__10076\,
            I => \N__10067\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10073\,
            I => \N__10064\
        );

    \I__2277\ : Span4Mux_v
    port map (
            O => \N__10070\,
            I => \N__10059\
        );

    \I__2276\ : LocalMux
    port map (
            O => \N__10067\,
            I => \N__10059\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__10064\,
            I => \N__10056\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__10059\,
            I => \N__10053\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__10056\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__2272\ : Odrv4
    port map (
            O => \N__10053\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__2271\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10045\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10042\
        );

    \I__2269\ : Span4Mux_v
    port map (
            O => \N__10042\,
            I => \N__10039\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__10039\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0\
        );

    \I__2267\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10031\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10035\,
            I => \N__10028\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__10034\,
            I => \N__10025\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__10022\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__10028\,
            I => \N__10019\
        );

    \I__2262\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10016\
        );

    \I__2261\ : Span4Mux_h
    port map (
            O => \N__10022\,
            I => \N__10011\
        );

    \I__2260\ : Span4Mux_v
    port map (
            O => \N__10019\,
            I => \N__10008\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10005\
        );

    \I__2258\ : InMux
    port map (
            O => \N__10015\,
            I => \N__10002\
        );

    \I__2257\ : InMux
    port map (
            O => \N__10014\,
            I => \N__9999\
        );

    \I__2256\ : Odrv4
    port map (
            O => \N__10011\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_EN\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__10008\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_EN\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__10005\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_EN\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__10002\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_EN\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9999\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_EN\
        );

    \I__2251\ : IoInMux
    port map (
            O => \N__9988\,
            I => \N__9985\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__9985\,
            I => \N__9982\
        );

    \I__2249\ : Span12Mux_s10_h
    port map (
            O => \N__9982\,
            I => \N__9979\
        );

    \I__2248\ : Odrv12
    port map (
            O => \N__9979\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__9976\,
            I => \U409_CIA.CLK_CIA6_4_cascade_\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__9973\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9966\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9963\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9957\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__9963\,
            I => \N__9957\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9962\,
            I => \N__9954\
        );

    \I__2240\ : Odrv12
    port map (
            O => \N__9957\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9954\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9944\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9941\
        );

    \I__2236\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9938\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9935\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__9941\,
            I => \N__9930\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9930\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__9935\,
            I => \N__9926\
        );

    \I__2231\ : Span4Mux_v
    port map (
            O => \N__9930\,
            I => \N__9923\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9929\,
            I => \N__9920\
        );

    \I__2229\ : Span4Mux_h
    port map (
            O => \N__9926\,
            I => \N__9916\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__9923\,
            I => \N__9911\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__9920\,
            I => \N__9911\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9908\
        );

    \I__2225\ : Odrv4
    port map (
            O => \N__9916\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2224\ : Odrv4
    port map (
            O => \N__9911\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9908\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__9898\,
            I => \N__9893\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9897\,
            I => \N__9890\
        );

    \I__2219\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9887\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__9893\,
            I => \N__9884\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9890\,
            I => \N__9879\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9887\,
            I => \N__9879\
        );

    \I__2215\ : Odrv4
    port map (
            O => \N__9884\,
            I => \CIA_SPACE\
        );

    \I__2214\ : Odrv12
    port map (
            O => \N__9879\,
            I => \CIA_SPACE\
        );

    \I__2213\ : IoInMux
    port map (
            O => \N__9874\,
            I => \N__9870\
        );

    \I__2212\ : IoInMux
    port map (
            O => \N__9873\,
            I => \N__9867\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__9870\,
            I => \N__9862\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9862\
        );

    \I__2209\ : IoSpan4Mux
    port map (
            O => \N__9862\,
            I => \N__9859\
        );

    \I__2208\ : Span4Mux_s2_v
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__9856\,
            I => \N__9852\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9855\,
            I => \N__9849\
        );

    \I__2205\ : Sp12to4
    port map (
            O => \N__9852\,
            I => \N__9845\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9849\,
            I => \N__9842\
        );

    \I__2203\ : CascadeMux
    port map (
            O => \N__9848\,
            I => \N__9839\
        );

    \I__2202\ : Span12Mux_v
    port map (
            O => \N__9845\,
            I => \N__9836\
        );

    \I__2201\ : Span4Mux_v
    port map (
            O => \N__9842\,
            I => \N__9833\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9830\
        );

    \I__2199\ : Odrv12
    port map (
            O => \N__9836\,
            I => \TACK_EN\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__9833\,
            I => \TACK_EN\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9830\,
            I => \TACK_EN\
        );

    \I__2196\ : IoInMux
    port map (
            O => \N__9823\,
            I => \N__9820\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9820\,
            I => \N__9817\
        );

    \I__2194\ : Span4Mux_s3_v
    port map (
            O => \N__9817\,
            I => \N__9814\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__9814\,
            I => \N__9811\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__9811\,
            I => \N__9808\
        );

    \I__2191\ : Sp12to4
    port map (
            O => \N__9808\,
            I => \N__9805\
        );

    \I__2190\ : Span12Mux_v
    port map (
            O => \N__9805\,
            I => \N__9802\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__9802\,
            I => \TCIn_1_i\
        );

    \I__2188\ : IoInMux
    port map (
            O => \N__9799\,
            I => \N__9795\
        );

    \I__2187\ : IoInMux
    port map (
            O => \N__9798\,
            I => \N__9792\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9795\,
            I => \N__9787\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9787\
        );

    \I__2184\ : IoSpan4Mux
    port map (
            O => \N__9787\,
            I => \N__9782\
        );

    \I__2183\ : IoInMux
    port map (
            O => \N__9786\,
            I => \N__9779\
        );

    \I__2182\ : IoInMux
    port map (
            O => \N__9785\,
            I => \N__9776\
        );

    \I__2181\ : IoSpan4Mux
    port map (
            O => \N__9782\,
            I => \N__9773\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9768\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9768\
        );

    \I__2178\ : IoSpan4Mux
    port map (
            O => \N__9773\,
            I => \N__9763\
        );

    \I__2177\ : IoSpan4Mux
    port map (
            O => \N__9768\,
            I => \N__9763\
        );

    \I__2176\ : Span4Mux_s0_h
    port map (
            O => \N__9763\,
            I => \N__9760\
        );

    \I__2175\ : Span4Mux_h
    port map (
            O => \N__9760\,
            I => \N__9756\
        );

    \I__2174\ : IoInMux
    port map (
            O => \N__9759\,
            I => \N__9753\
        );

    \I__2173\ : Span4Mux_h
    port map (
            O => \N__9756\,
            I => \N__9750\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9753\,
            I => \N__9747\
        );

    \I__2171\ : Span4Mux_h
    port map (
            O => \N__9750\,
            I => \N__9742\
        );

    \I__2170\ : Span4Mux_s2_v
    port map (
            O => \N__9747\,
            I => \N__9742\
        );

    \I__2169\ : Span4Mux_v
    port map (
            O => \N__9742\,
            I => \N__9739\
        );

    \I__2168\ : Odrv4
    port map (
            O => \N__9739\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2167\ : SRMux
    port map (
            O => \N__9736\,
            I => \N__9703\
        );

    \I__2166\ : SRMux
    port map (
            O => \N__9735\,
            I => \N__9703\
        );

    \I__2165\ : SRMux
    port map (
            O => \N__9734\,
            I => \N__9703\
        );

    \I__2164\ : SRMux
    port map (
            O => \N__9733\,
            I => \N__9703\
        );

    \I__2163\ : SRMux
    port map (
            O => \N__9732\,
            I => \N__9703\
        );

    \I__2162\ : SRMux
    port map (
            O => \N__9731\,
            I => \N__9703\
        );

    \I__2161\ : SRMux
    port map (
            O => \N__9730\,
            I => \N__9703\
        );

    \I__2160\ : SRMux
    port map (
            O => \N__9729\,
            I => \N__9703\
        );

    \I__2159\ : SRMux
    port map (
            O => \N__9728\,
            I => \N__9703\
        );

    \I__2158\ : SRMux
    port map (
            O => \N__9727\,
            I => \N__9703\
        );

    \I__2157\ : SRMux
    port map (
            O => \N__9726\,
            I => \N__9703\
        );

    \I__2156\ : GlobalMux
    port map (
            O => \N__9703\,
            I => \N__9700\
        );

    \I__2155\ : gio2CtrlBuf
    port map (
            O => \N__9700\,
            I => \RESETn_c_i_g\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__9697\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9691\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__9691\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9684\
        );

    \I__2150\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9681\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9684\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9681\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9676\,
            I => \N__9670\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9675\,
            I => \N__9665\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9665\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9673\,
            I => \N__9662\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9670\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9665\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9662\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__9654\,
            I => \N__9646\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9641\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9641\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9649\,
            I => \N__9638\
        );

    \I__2135\ : InMux
    port map (
            O => \N__9646\,
            I => \N__9635\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__9641\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__9638\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9635\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__2131\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9624\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9627\,
            I => \N__9621\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9624\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__9621\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__9616\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__2126\ : IoInMux
    port map (
            O => \N__9613\,
            I => \N__9609\
        );

    \I__2125\ : IoInMux
    port map (
            O => \N__9612\,
            I => \N__9606\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9609\,
            I => \N__9601\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__9606\,
            I => \N__9601\
        );

    \I__2122\ : IoSpan4Mux
    port map (
            O => \N__9601\,
            I => \N__9597\
        );

    \I__2121\ : IoInMux
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__2120\ : Span4Mux_s3_v
    port map (
            O => \N__9597\,
            I => \N__9591\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__9594\,
            I => \N__9588\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__9591\,
            I => \N__9583\
        );

    \I__2117\ : Span4Mux_s3_v
    port map (
            O => \N__9588\,
            I => \N__9583\
        );

    \I__2116\ : Sp12to4
    port map (
            O => \N__9583\,
            I => \N__9580\
        );

    \I__2115\ : Span12Mux_h
    port map (
            O => \N__9580\,
            I => \N__9577\
        );

    \I__2114\ : Span12Mux_v
    port map (
            O => \N__9577\,
            I => \N__9572\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9567\
        );

    \I__2112\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9567\
        );

    \I__2111\ : Odrv12
    port map (
            O => \N__9572\,
            I => \TACK_OUTn\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9567\,
            I => \TACK_OUTn\
        );

    \I__2109\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9558\
        );

    \I__2108\ : InMux
    port map (
            O => \N__9561\,
            I => \N__9555\
        );

    \I__2107\ : LocalMux
    port map (
            O => \N__9558\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__9555\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__2105\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9545\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9540\
        );

    \I__2103\ : InMux
    port map (
            O => \N__9548\,
            I => \N__9540\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__9545\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9540\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9532\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9532\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__2098\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9524\
        );

    \I__2097\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9521\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9518\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__9524\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9521\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9518\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9511\,
            I => \N__9507\
        );

    \I__2091\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9504\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9507\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9504\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9499\,
            I => \N__9494\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9489\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9485\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9494\,
            I => \N__9482\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9493\,
            I => \N__9479\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9476\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9472\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9469\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9485\,
            I => \N__9466\
        );

    \I__2079\ : Span4Mux_v
    port map (
            O => \N__9482\,
            I => \N__9461\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9479\,
            I => \N__9461\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9476\,
            I => \N__9458\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9475\,
            I => \N__9455\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__9472\,
            I => \N__9450\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9469\,
            I => \N__9450\
        );

    \I__2073\ : Span4Mux_v
    port map (
            O => \N__9466\,
            I => \N__9447\
        );

    \I__2072\ : Span4Mux_h
    port map (
            O => \N__9461\,
            I => \N__9440\
        );

    \I__2071\ : Span4Mux_v
    port map (
            O => \N__9458\,
            I => \N__9440\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9455\,
            I => \N__9440\
        );

    \I__2069\ : Span4Mux_v
    port map (
            O => \N__9450\,
            I => \N__9437\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__9447\,
            I => \N__9432\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__9440\,
            I => \N__9432\
        );

    \I__2066\ : Sp12to4
    port map (
            O => \N__9437\,
            I => \N__9427\
        );

    \I__2065\ : Sp12to4
    port map (
            O => \N__9432\,
            I => \N__9427\
        );

    \I__2064\ : Span12Mux_h
    port map (
            O => \N__9427\,
            I => \N__9424\
        );

    \I__2063\ : Span12Mux_v
    port map (
            O => \N__9424\,
            I => \N__9421\
        );

    \I__2062\ : Odrv12
    port map (
            O => \N__9421\,
            I => \TSn_c\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9418\,
            I => \N__9401\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9417\,
            I => \N__9401\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9401\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9401\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9401\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9413\,
            I => \N__9396\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9412\,
            I => \N__9396\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__9401\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9396\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9388\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__9388\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9385\,
            I => \N__9382\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9376\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__2046\ : Sp12to4
    port map (
            O => \N__9373\,
            I => \N__9370\
        );

    \I__2045\ : Span12Mux_h
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__2044\ : Span12Mux_v
    port map (
            O => \N__9367\,
            I => \N__9364\
        );

    \I__2043\ : Odrv12
    port map (
            O => \N__9364\,
            I => \TACKn_in\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__9361\,
            I => \N__9358\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9355\,
            I => \N__9351\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9354\,
            I => \N__9348\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__9351\,
            I => \N__9343\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__9348\,
            I => \N__9343\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__9343\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__2035\ : IoInMux
    port map (
            O => \N__9340\,
            I => \N__9337\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__2033\ : Span12Mux_s1_v
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__2032\ : Span12Mux_h
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__2031\ : Odrv12
    port map (
            O => \N__9328\,
            I => \BUFENn_c\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9319\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9319\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__2027\ : Span4Mux_v
    port map (
            O => \N__9316\,
            I => \N__9312\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9309\
        );

    \I__2025\ : Odrv4
    port map (
            O => \N__9312\,
            I => \U409_ADDRESS_DECODE_un2_REGSPACEn_0\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__9309\,
            I => \U409_ADDRESS_DECODE_un2_REGSPACEn_0\
        );

    \I__2023\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9298\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9298\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9298\,
            I => \N__9292\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9286\
        );

    \I__2019\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9286\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9283\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__9292\,
            I => \N__9280\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9291\,
            I => \N__9277\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9286\,
            I => \N__9271\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9271\
        );

    \I__2013\ : Span4Mux_v
    port map (
            O => \N__9280\,
            I => \N__9266\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__9277\,
            I => \N__9266\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9276\,
            I => \N__9263\
        );

    \I__2010\ : Span4Mux_v
    port map (
            O => \N__9271\,
            I => \N__9260\
        );

    \I__2009\ : Span4Mux_h
    port map (
            O => \N__9266\,
            I => \N__9257\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9263\,
            I => \N__9254\
        );

    \I__2007\ : Sp12to4
    port map (
            O => \N__9260\,
            I => \N__9251\
        );

    \I__2006\ : Span4Mux_v
    port map (
            O => \N__9257\,
            I => \N__9248\
        );

    \I__2005\ : Span4Mux_v
    port map (
            O => \N__9254\,
            I => \N__9245\
        );

    \I__2004\ : Odrv12
    port map (
            O => \N__9251\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__9248\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__9245\,
            I => \U409_ADDRESS_DECODE_Z2_SPACE\
        );

    \I__2001\ : IoInMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__1999\ : IoSpan4Mux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__1998\ : Sp12to4
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__1997\ : Span12Mux_v
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__9223\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9220\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__1994\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9211\
        );

    \I__1992\ : Span4Mux_v
    port map (
            O => \N__9211\,
            I => \N__9208\
        );

    \I__1991\ : Sp12to4
    port map (
            O => \N__9208\,
            I => \N__9205\
        );

    \I__1990\ : Span12Mux_h
    port map (
            O => \N__9205\,
            I => \N__9202\
        );

    \I__1989\ : Odrv12
    port map (
            O => \N__9202\,
            I => \A_c_12\
        );

    \I__1988\ : IoInMux
    port map (
            O => \N__9199\,
            I => \N__9196\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__1986\ : Span4Mux_s1_h
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__1985\ : Sp12to4
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__1984\ : Span12Mux_s8_v
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1983\ : Span12Mux_h
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__1982\ : Odrv12
    port map (
            O => \N__9181\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__9175\,
            I => \CIA_ENABLE\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1977\ : Span4Mux_v
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__1976\ : Sp12to4
    port map (
            O => \N__9163\,
            I => \N__9160\
        );

    \I__1975\ : Span12Mux_h
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__1974\ : Odrv12
    port map (
            O => \N__9157\,
            I => \A_c_13\
        );

    \I__1973\ : IoInMux
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__1971\ : IoSpan4Mux
    port map (
            O => \N__9148\,
            I => \N__9145\
        );

    \I__1970\ : IoSpan4Mux
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__1969\ : Sp12to4
    port map (
            O => \N__9142\,
            I => \N__9139\
        );

    \I__1968\ : Span12Mux_s7_h
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__1967\ : Odrv12
    port map (
            O => \N__9136\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__9133\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__9130\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__1963\ : InMux
    port map (
            O => \N__9126\,
            I => \N__9116\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9116\
        );

    \I__1961\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9111\
        );

    \I__1960\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9111\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__9116\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__9111\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1957\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9100\
        );

    \I__1956\ : InMux
    port map (
            O => \N__9105\,
            I => \N__9100\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__9100\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__9097\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__1953\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9079\
        );

    \I__1952\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9079\
        );

    \I__1951\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9079\
        );

    \I__1950\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9079\
        );

    \I__1949\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9079\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__9079\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__9076\,
            I => \N__9071\
        );

    \I__1946\ : CascadeMux
    port map (
            O => \N__9075\,
            I => \N__9068\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__9074\,
            I => \N__9065\
        );

    \I__1944\ : InMux
    port map (
            O => \N__9071\,
            I => \N__9055\
        );

    \I__1943\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9055\
        );

    \I__1942\ : InMux
    port map (
            O => \N__9065\,
            I => \N__9055\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9055\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__9055\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__9052\,
            I => \N__9047\
        );

    \I__1938\ : InMux
    port map (
            O => \N__9051\,
            I => \N__9041\
        );

    \I__1937\ : InMux
    port map (
            O => \N__9050\,
            I => \N__9041\
        );

    \I__1936\ : InMux
    port map (
            O => \N__9047\,
            I => \N__9038\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9035\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__9041\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__9038\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__9035\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__9028\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9019\
        );

    \I__1929\ : InMux
    port map (
            O => \N__9024\,
            I => \N__9016\
        );

    \I__1928\ : InMux
    port map (
            O => \N__9023\,
            I => \N__9011\
        );

    \I__1927\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9011\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__9019\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__9016\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__9011\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1923\ : InMux
    port map (
            O => \N__9004\,
            I => \N__8998\
        );

    \I__1922\ : InMux
    port map (
            O => \N__9003\,
            I => \N__8998\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__8995\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__8992\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8982\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8982\
        );

    \I__1916\ : InMux
    port map (
            O => \N__8987\,
            I => \N__8979\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8982\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8979\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__8974\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8968\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8968\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8959\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8959\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1907\ : InMux
    port map (
            O => \N__8956\,
            I => \N__8953\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8953\,
            I => \N__8949\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8952\,
            I => \N__8946\
        );

    \I__1904\ : Span4Mux_v
    port map (
            O => \N__8949\,
            I => \N__8941\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8946\,
            I => \N__8941\
        );

    \I__1902\ : Span4Mux_v
    port map (
            O => \N__8941\,
            I => \N__8937\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8934\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__8937\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__8934\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__8929\,
            I => \N__8926\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8922\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8925\,
            I => \N__8919\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8922\,
            I => \N__8914\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8914\
        );

    \I__1893\ : Span4Mux_h
    port map (
            O => \N__8914\,
            I => \N__8911\
        );

    \I__1892\ : Span4Mux_v
    port map (
            O => \N__8911\,
            I => \N__8908\
        );

    \I__1891\ : Span4Mux_v
    port map (
            O => \N__8908\,
            I => \N__8905\
        );

    \I__1890\ : Odrv4
    port map (
            O => \N__8905\,
            I => \AUTOVECTOR\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8899\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8899\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8893\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8893\,
            I => \N__8890\
        );

    \I__1885\ : Span4Mux_h
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1884\ : Span4Mux_h
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__1883\ : Odrv4
    port map (
            O => \N__8884\,
            I => \AC_TACK\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__8881\,
            I => \N__8878\
        );

    \I__1881\ : InMux
    port map (
            O => \N__8878\,
            I => \N__8874\
        );

    \I__1880\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8871\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8874\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8871\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__8866\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__8863\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8856\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8859\,
            I => \N__8853\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8850\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8853\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8850\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1870\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8842\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8842\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8836\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8836\,
            I => \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d\
        );

    \I__1866\ : IoInMux
    port map (
            O => \N__8833\,
            I => \N__8830\
        );

    \I__1865\ : LocalMux
    port map (
            O => \N__8830\,
            I => \N__8827\
        );

    \I__1864\ : IoSpan4Mux
    port map (
            O => \N__8827\,
            I => \N__8824\
        );

    \I__1863\ : Sp12to4
    port map (
            O => \N__8824\,
            I => \N__8821\
        );

    \I__1862\ : Span12Mux_s6_v
    port map (
            O => \N__8821\,
            I => \N__8818\
        );

    \I__1861\ : Span12Mux_v
    port map (
            O => \N__8818\,
            I => \N__8814\
        );

    \I__1860\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8811\
        );

    \I__1859\ : Odrv12
    port map (
            O => \N__8814\,
            I => \ROMENn_c\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__8811\,
            I => \ROMENn_c\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__8806\,
            I => \N__8803\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8803\,
            I => \N__8799\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8802\,
            I => \N__8796\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8799\,
            I => \N__8790\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8783\
        );

    \I__1851\ : Span4Mux_h
    port map (
            O => \N__8790\,
            I => \N__8780\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8789\,
            I => \N__8777\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8788\,
            I => \N__8770\
        );

    \I__1848\ : InMux
    port map (
            O => \N__8787\,
            I => \N__8770\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8770\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__8783\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__8780\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1844\ : LocalMux
    port map (
            O => \N__8777\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__8770\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8758\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8758\,
            I => \N__8755\
        );

    \I__1840\ : Span4Mux_h
    port map (
            O => \N__8755\,
            I => \N__8746\
        );

    \I__1839\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8743\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8740\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8752\,
            I => \N__8737\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8730\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8730\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8749\,
            I => \N__8730\
        );

    \I__1833\ : Odrv4
    port map (
            O => \N__8746\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8743\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8740\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8737\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8730\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__8719\,
            I => \N__8716\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8716\,
            I => \N__8713\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8713\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8706\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8709\,
            I => \N__8703\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__8706\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8703\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8695\,
            I => \N__8692\
        );

    \I__1819\ : Odrv4
    port map (
            O => \N__8692\,
            I => \U409_TRANSFER_ACK.G_14_0_o7_6\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__8689\,
            I => \U409_TRANSFER_ACK.G_14_0_4_cascade_\
        );

    \I__1817\ : InMux
    port map (
            O => \N__8686\,
            I => \N__8683\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8683\,
            I => \U409_TRANSFER_ACK.g0_0_0_o6_4\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__8680\,
            I => \N__8677\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8671\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8671\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8671\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8668\,
            I => \N__8664\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__8667\,
            I => \N__8658\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8653\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8650\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8641\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8641\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8641\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8641\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8638\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8653\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8650\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8641\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8638\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__8629\,
            I => \N__8620\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__8628\,
            I => \N__8617\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8614\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8611\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8602\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8624\,
            I => \N__8602\
        );

    \I__1792\ : InMux
    port map (
            O => \N__8623\,
            I => \N__8602\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8602\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8617\,
            I => \N__8599\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8614\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__8611\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8602\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8599\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8585\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8580\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8580\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8585\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8580\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__1780\ : CascadeMux
    port map (
            O => \N__8575\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8567\
        );

    \I__1778\ : InMux
    port map (
            O => \N__8571\,
            I => \N__8564\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8561\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__8567\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__8564\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__8561\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8554\,
            I => \N__8551\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8551\,
            I => \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8539\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8547\,
            I => \N__8533\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8528\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8545\,
            I => \N__8523\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8523\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8517\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8517\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8539\,
            I => \N__8514\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8538\,
            I => \N__8509\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8509\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8506\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8502\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8497\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8497\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8492\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8523\,
            I => \N__8492\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8522\,
            I => \N__8489\
        );

    \I__1754\ : LocalMux
    port map (
            O => \N__8517\,
            I => \N__8485\
        );

    \I__1753\ : Span4Mux_h
    port map (
            O => \N__8514\,
            I => \N__8478\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8478\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8478\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8475\
        );

    \I__1749\ : Span4Mux_v
    port map (
            O => \N__8502\,
            I => \N__8466\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8466\
        );

    \I__1747\ : Span4Mux_v
    port map (
            O => \N__8492\,
            I => \N__8466\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8466\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8463\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__8485\,
            I => \N__8460\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__8478\,
            I => \N__8455\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8455\
        );

    \I__1741\ : Span4Mux_h
    port map (
            O => \N__8466\,
            I => \N__8450\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__8463\,
            I => \N__8450\
        );

    \I__1739\ : Span4Mux_v
    port map (
            O => \N__8460\,
            I => \N__8445\
        );

    \I__1738\ : Span4Mux_v
    port map (
            O => \N__8455\,
            I => \N__8445\
        );

    \I__1737\ : Span4Mux_v
    port map (
            O => \N__8450\,
            I => \N__8442\
        );

    \I__1736\ : Sp12to4
    port map (
            O => \N__8445\,
            I => \N__8437\
        );

    \I__1735\ : Sp12to4
    port map (
            O => \N__8442\,
            I => \N__8437\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8437\,
            I => \A_c_21\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8430\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8427\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8421\
        );

    \I__1729\ : Span4Mux_v
    port map (
            O => \N__8424\,
            I => \N__8413\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__8421\,
            I => \N__8413\
        );

    \I__1727\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8410\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8419\,
            I => \N__8407\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8404\
        );

    \I__1724\ : Sp12to4
    port map (
            O => \N__8413\,
            I => \N__8399\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8410\,
            I => \N__8399\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8407\,
            I => \N__8394\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8404\,
            I => \N__8394\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__8399\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1719\ : Odrv4
    port map (
            O => \N__8394\,
            I => \U409_ADDRESS_DECODE_ROMEN_1\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8384\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8388\,
            I => \N__8381\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__8387\,
            I => \N__8378\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__8384\,
            I => \N__8374\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__8381\,
            I => \N__8371\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8368\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \N__8365\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8374\,
            I => \N__8362\
        );

    \I__1710\ : Span4Mux_h
    port map (
            O => \N__8371\,
            I => \N__8359\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8356\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8353\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__8362\,
            I => \N__8350\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__8359\,
            I => \N__8347\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__8356\,
            I => \N__8344\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8353\,
            I => \N__8341\
        );

    \I__1703\ : Sp12to4
    port map (
            O => \N__8350\,
            I => \N__8338\
        );

    \I__1702\ : Sp12to4
    port map (
            O => \N__8347\,
            I => \N__8333\
        );

    \I__1701\ : Sp12to4
    port map (
            O => \N__8344\,
            I => \N__8333\
        );

    \I__1700\ : Span12Mux_h
    port map (
            O => \N__8341\,
            I => \N__8330\
        );

    \I__1699\ : Span12Mux_h
    port map (
            O => \N__8338\,
            I => \N__8327\
        );

    \I__1698\ : Span12Mux_v
    port map (
            O => \N__8333\,
            I => \N__8324\
        );

    \I__1697\ : Span12Mux_v
    port map (
            O => \N__8330\,
            I => \N__8321\
        );

    \I__1696\ : Span12Mux_v
    port map (
            O => \N__8327\,
            I => \N__8316\
        );

    \I__1695\ : Span12Mux_h
    port map (
            O => \N__8324\,
            I => \N__8316\
        );

    \I__1694\ : Odrv12
    port map (
            O => \N__8321\,
            I => \OVL_c\
        );

    \I__1693\ : Odrv12
    port map (
            O => \N__8316\,
            I => \OVL_c\
        );

    \I__1692\ : InMux
    port map (
            O => \N__8311\,
            I => \N__8308\
        );

    \I__1691\ : LocalMux
    port map (
            O => \N__8308\,
            I => \N__8305\
        );

    \I__1690\ : Span12Mux_v
    port map (
            O => \N__8305\,
            I => \N__8301\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8304\,
            I => \N__8298\
        );

    \I__1688\ : Odrv12
    port map (
            O => \N__8301\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8298\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\
        );

    \I__1686\ : CascadeMux
    port map (
            O => \N__8293\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_\
        );

    \I__1685\ : IoInMux
    port map (
            O => \N__8290\,
            I => \N__8287\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8287\,
            I => \N__8284\
        );

    \I__1683\ : IoSpan4Mux
    port map (
            O => \N__8284\,
            I => \N__8281\
        );

    \I__1682\ : IoSpan4Mux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1681\ : Span4Mux_s1_v
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1680\ : Sp12to4
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8272\,
            I => \PORTSIZE_0_i\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8269\,
            I => \U409_TRANSFER_ACK.G_14_0_o7_2_cascade_\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8263\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__8260\,
            I => \N__8257\
        );

    \I__1674\ : Odrv4
    port map (
            O => \N__8257\,
            I => \U409_TRANSFER_ACK.G_14_0_o7_4\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__8253\,
            I => \N__8245\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__8252\,
            I => \N__8242\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8238\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__8248\,
            I => \N__8233\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8230\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8227\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__8241\,
            I => \N__8224\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__8238\,
            I => \N__8218\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__8237\,
            I => \N__8212\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__8236\,
            I => \N__8209\
        );

    \I__1662\ : Span4Mux_h
    port map (
            O => \N__8233\,
            I => \N__8202\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__8230\,
            I => \N__8202\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8227\,
            I => \N__8202\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8199\
        );

    \I__1658\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8194\
        );

    \I__1657\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8194\
        );

    \I__1656\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8191\
        );

    \I__1655\ : Span4Mux_v
    port map (
            O => \N__8218\,
            I => \N__8188\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8217\,
            I => \N__8183\
        );

    \I__1653\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8183\
        );

    \I__1652\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8180\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8177\
        );

    \I__1650\ : InMux
    port map (
            O => \N__8209\,
            I => \N__8174\
        );

    \I__1649\ : Span4Mux_v
    port map (
            O => \N__8202\,
            I => \N__8167\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8167\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8194\,
            I => \N__8167\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__8191\,
            I => \N__8164\
        );

    \I__1645\ : Span4Mux_v
    port map (
            O => \N__8188\,
            I => \N__8159\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__8183\,
            I => \N__8159\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__8180\,
            I => \N__8156\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8153\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__8174\,
            I => \N__8150\
        );

    \I__1640\ : Span4Mux_v
    port map (
            O => \N__8167\,
            I => \N__8145\
        );

    \I__1639\ : Span4Mux_v
    port map (
            O => \N__8164\,
            I => \N__8145\
        );

    \I__1638\ : Span4Mux_h
    port map (
            O => \N__8159\,
            I => \N__8138\
        );

    \I__1637\ : Span4Mux_v
    port map (
            O => \N__8156\,
            I => \N__8138\
        );

    \I__1636\ : Span4Mux_v
    port map (
            O => \N__8153\,
            I => \N__8138\
        );

    \I__1635\ : Span12Mux_v
    port map (
            O => \N__8150\,
            I => \N__8131\
        );

    \I__1634\ : Sp12to4
    port map (
            O => \N__8145\,
            I => \N__8131\
        );

    \I__1633\ : Sp12to4
    port map (
            O => \N__8138\,
            I => \N__8131\
        );

    \I__1632\ : Odrv12
    port map (
            O => \N__8131\,
            I => \A_c_20\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8128\,
            I => \N__8123\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__8127\,
            I => \N__8120\
        );

    \I__1629\ : InMux
    port map (
            O => \N__8126\,
            I => \N__8116\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8123\,
            I => \N__8113\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8110\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8119\,
            I => \N__8107\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8116\,
            I => \ATA_BASE_7\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8113\,
            I => \ATA_BASE_7\
        );

    \I__1623\ : LocalMux
    port map (
            O => \N__8110\,
            I => \ATA_BASE_7\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__8107\,
            I => \ATA_BASE_7\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8093\
        );

    \I__1620\ : InMux
    port map (
            O => \N__8097\,
            I => \N__8089\
        );

    \I__1619\ : InMux
    port map (
            O => \N__8096\,
            I => \N__8086\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8083\
        );

    \I__1617\ : InMux
    port map (
            O => \N__8092\,
            I => \N__8080\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__8089\,
            I => \N__8077\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__8086\,
            I => \ATA_BASE_4\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__8083\,
            I => \ATA_BASE_4\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__8080\,
            I => \ATA_BASE_4\
        );

    \I__1612\ : Odrv4
    port map (
            O => \N__8077\,
            I => \ATA_BASE_4\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8068\,
            I => \N__8065\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__8065\,
            I => \U409_TRANSFER_ACK.G_14_0_o7_3\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__8059\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0\
        );

    \I__1607\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8052\
        );

    \I__1606\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8049\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8052\,
            I => \U409_TRANSFER_ACK.N_13\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__8049\,
            I => \U409_TRANSFER_ACK.N_13\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__8044\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8037\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__8040\,
            I => \N__8034\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__8037\,
            I => \N__8025\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8022\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8019\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8014\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8031\,
            I => \N__8011\
        );

    \I__1595\ : InMux
    port map (
            O => \N__8030\,
            I => \N__8005\
        );

    \I__1594\ : InMux
    port map (
            O => \N__8029\,
            I => \N__8005\
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__8028\,
            I => \N__8001\
        );

    \I__1592\ : Span4Mux_h
    port map (
            O => \N__8025\,
            I => \N__7994\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__8022\,
            I => \N__7994\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__8019\,
            I => \N__7994\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8018\,
            I => \N__7991\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8017\,
            I => \N__7988\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7983\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__7983\
        );

    \I__1585\ : InMux
    port map (
            O => \N__8010\,
            I => \N__7980\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__7977\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7974\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7970\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__7994\,
            I => \N__7964\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7964\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7988\,
            I => \N__7961\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__7983\,
            I => \N__7952\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7980\,
            I => \N__7952\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__7977\,
            I => \N__7952\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7974\,
            I => \N__7952\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7973\,
            I => \N__7949\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__7970\,
            I => \N__7946\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7943\
        );

    \I__1571\ : Span4Mux_v
    port map (
            O => \N__7964\,
            I => \N__7940\
        );

    \I__1570\ : Span4Mux_v
    port map (
            O => \N__7961\,
            I => \N__7933\
        );

    \I__1569\ : Span4Mux_h
    port map (
            O => \N__7952\,
            I => \N__7933\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7949\,
            I => \N__7933\
        );

    \I__1567\ : Sp12to4
    port map (
            O => \N__7946\,
            I => \N__7928\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7928\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__7940\,
            I => \N__7925\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__7933\,
            I => \N__7922\
        );

    \I__1563\ : Span12Mux_v
    port map (
            O => \N__7928\,
            I => \N__7919\
        );

    \I__1562\ : Sp12to4
    port map (
            O => \N__7925\,
            I => \N__7914\
        );

    \I__1561\ : Sp12to4
    port map (
            O => \N__7922\,
            I => \N__7914\
        );

    \I__1560\ : Odrv12
    port map (
            O => \N__7919\,
            I => \A_c_23\
        );

    \I__1559\ : Odrv12
    port map (
            O => \N__7914\,
            I => \A_c_23\
        );

    \I__1558\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7906\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7906\,
            I => \N__7903\
        );

    \I__1556\ : Odrv4
    port map (
            O => \N__7903\,
            I => \U409_TRANSFER_ACK.N_24\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__7900\,
            I => \N__7897\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__7888\,
            I => \U409_TRANSFER_ACK.G_14_0_1_1\
        );

    \I__1550\ : CascadeMux
    port map (
            O => \N__7885\,
            I => \U409_TRANSFER_ACK.G_14_0_1_cascade_\
        );

    \I__1549\ : CascadeMux
    port map (
            O => \N__7882\,
            I => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7879\,
            I => \N__7871\
        );

    \I__1547\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7871\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__7877\,
            I => \N__7866\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7863\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__7871\,
            I => \N__7859\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__7870\,
            I => \N__7856\
        );

    \I__1542\ : InMux
    port map (
            O => \N__7869\,
            I => \N__7851\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7866\,
            I => \N__7851\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7863\,
            I => \N__7848\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7862\,
            I => \N__7845\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__7859\,
            I => \N__7842\
        );

    \I__1537\ : InMux
    port map (
            O => \N__7856\,
            I => \N__7839\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__7851\,
            I => \N__7835\
        );

    \I__1535\ : Span4Mux_v
    port map (
            O => \N__7848\,
            I => \N__7830\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__7845\,
            I => \N__7830\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__7842\,
            I => \N__7825\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__7839\,
            I => \N__7825\
        );

    \I__1531\ : InMux
    port map (
            O => \N__7838\,
            I => \N__7819\
        );

    \I__1530\ : Span4Mux_v
    port map (
            O => \N__7835\,
            I => \N__7816\
        );

    \I__1529\ : Span4Mux_v
    port map (
            O => \N__7830\,
            I => \N__7813\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__7825\,
            I => \N__7810\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7824\,
            I => \N__7805\
        );

    \I__1526\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7805\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7802\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7819\,
            I => \N__7789\
        );

    \I__1523\ : Sp12to4
    port map (
            O => \N__7816\,
            I => \N__7789\
        );

    \I__1522\ : Sp12to4
    port map (
            O => \N__7813\,
            I => \N__7789\
        );

    \I__1521\ : Sp12to4
    port map (
            O => \N__7810\,
            I => \N__7789\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7805\,
            I => \N__7789\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7789\
        );

    \I__1518\ : Span12Mux_h
    port map (
            O => \N__7789\,
            I => \N__7786\
        );

    \I__1517\ : Span12Mux_v
    port map (
            O => \N__7786\,
            I => \N__7783\
        );

    \I__1516\ : Odrv12
    port map (
            O => \N__7783\,
            I => \A_c_19\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__7779\,
            I => \N__7771\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__7778\,
            I => \N__7767\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__7777\,
            I => \N__7764\
        );

    \I__1511\ : InMux
    port map (
            O => \N__7774\,
            I => \N__7761\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7771\,
            I => \N__7758\
        );

    \I__1509\ : InMux
    port map (
            O => \N__7770\,
            I => \N__7755\
        );

    \I__1508\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7750\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7750\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7761\,
            I => \N__7747\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__7758\,
            I => \N__7742\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__7755\,
            I => \N__7742\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7750\,
            I => \N__7739\
        );

    \I__1502\ : Span4Mux_v
    port map (
            O => \N__7747\,
            I => \N__7736\
        );

    \I__1501\ : Span4Mux_v
    port map (
            O => \N__7742\,
            I => \N__7731\
        );

    \I__1500\ : Span12Mux_v
    port map (
            O => \N__7739\,
            I => \N__7726\
        );

    \I__1499\ : Sp12to4
    port map (
            O => \N__7736\,
            I => \N__7726\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7723\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7720\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7731\,
            I => \N__7717\
        );

    \I__1495\ : Span12Mux_s11_h
    port map (
            O => \N__7726\,
            I => \N__7710\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7710\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7720\,
            I => \N__7710\
        );

    \I__1492\ : Span4Mux_v
    port map (
            O => \N__7717\,
            I => \N__7707\
        );

    \I__1491\ : Span12Mux_v
    port map (
            O => \N__7710\,
            I => \N__7702\
        );

    \I__1490\ : Sp12to4
    port map (
            O => \N__7707\,
            I => \N__7702\
        );

    \I__1489\ : Odrv12
    port map (
            O => \N__7702\,
            I => \A_c_18\
        );

    \I__1488\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7696\,
            I => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7690\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7690\,
            I => \U409_ADDRESS_DECODE.REG_SPACE_3\
        );

    \I__1484\ : InMux
    port map (
            O => \N__7687\,
            I => \N__7684\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__7684\,
            I => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\
        );

    \I__1482\ : IoInMux
    port map (
            O => \N__7681\,
            I => \N__7678\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7678\,
            I => \N__7675\
        );

    \I__1480\ : Span12Mux_s0_v
    port map (
            O => \N__7675\,
            I => \N__7672\
        );

    \I__1479\ : Span12Mux_v
    port map (
            O => \N__7672\,
            I => \N__7669\
        );

    \I__1478\ : Odrv12
    port map (
            O => \N__7669\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7666\,
            I => \N__7662\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__7665\,
            I => \N__7655\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__7662\,
            I => \N__7651\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7661\,
            I => \N__7648\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7660\,
            I => \N__7645\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7659\,
            I => \N__7640\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7640\
        );

    \I__1470\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7635\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7635\
        );

    \I__1468\ : Span4Mux_h
    port map (
            O => \N__7651\,
            I => \N__7630\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__7648\,
            I => \N__7630\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7645\,
            I => \N__7625\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__7640\,
            I => \N__7625\
        );

    \I__1464\ : LocalMux
    port map (
            O => \N__7635\,
            I => \N__7622\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__7630\,
            I => \N__7616\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__7625\,
            I => \N__7616\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__7622\,
            I => \N__7613\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7610\
        );

    \I__1459\ : Sp12to4
    port map (
            O => \N__7616\,
            I => \N__7603\
        );

    \I__1458\ : Sp12to4
    port map (
            O => \N__7613\,
            I => \N__7603\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7610\,
            I => \N__7603\
        );

    \I__1456\ : Span12Mux_v
    port map (
            O => \N__7603\,
            I => \N__7600\
        );

    \I__1455\ : Odrv12
    port map (
            O => \N__7600\,
            I => \A_c_17\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__7597\,
            I => \N__7592\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__7596\,
            I => \N__7589\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7595\,
            I => \N__7585\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7592\,
            I => \N__7582\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7577\
        );

    \I__1449\ : InMux
    port map (
            O => \N__7588\,
            I => \N__7577\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7585\,
            I => \ATA_BASE_1\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7582\,
            I => \ATA_BASE_1\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7577\,
            I => \ATA_BASE_1\
        );

    \I__1445\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7566\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7569\,
            I => \N__7563\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7566\,
            I => \U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__7563\,
            I => \U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__7558\,
            I => \N__7553\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7557\,
            I => \N__7549\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7556\,
            I => \N__7546\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7553\,
            I => \N__7541\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7552\,
            I => \N__7541\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7549\,
            I => \N__7537\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7546\,
            I => \N__7534\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7531\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7528\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__7537\,
            I => \N__7525\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__7534\,
            I => \N__7522\
        );

    \I__1430\ : Span4Mux_v
    port map (
            O => \N__7531\,
            I => \N__7517\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7528\,
            I => \N__7517\
        );

    \I__1428\ : Sp12to4
    port map (
            O => \N__7525\,
            I => \N__7512\
        );

    \I__1427\ : Sp12to4
    port map (
            O => \N__7522\,
            I => \N__7512\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__7517\,
            I => \N__7509\
        );

    \I__1425\ : Span12Mux_h
    port map (
            O => \N__7512\,
            I => \N__7506\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__7509\,
            I => \N__7503\
        );

    \I__1423\ : Span12Mux_v
    port map (
            O => \N__7506\,
            I => \N__7500\
        );

    \I__1422\ : Sp12to4
    port map (
            O => \N__7503\,
            I => \N__7497\
        );

    \I__1421\ : Odrv12
    port map (
            O => \N__7500\,
            I => \A_c_16\
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__7497\,
            I => \A_c_16\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7492\,
            I => \N__7483\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7491\,
            I => \N__7478\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7490\,
            I => \N__7475\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7489\,
            I => \N__7472\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7488\,
            I => \N__7469\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7487\,
            I => \N__7466\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7486\,
            I => \N__7463\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7483\,
            I => \N__7458\
        );

    \I__1411\ : InMux
    port map (
            O => \N__7482\,
            I => \N__7455\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7452\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__7478\,
            I => \N__7445\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7475\,
            I => \N__7445\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7472\,
            I => \N__7442\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7469\,
            I => \N__7439\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7466\,
            I => \N__7436\
        );

    \I__1404\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7433\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7462\,
            I => \N__7428\
        );

    \I__1402\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7428\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__7458\,
            I => \N__7421\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7455\,
            I => \N__7421\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7421\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7418\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7415\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__7445\,
            I => \N__7411\
        );

    \I__1395\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7406\
        );

    \I__1394\ : Span4Mux_v
    port map (
            O => \N__7439\,
            I => \N__7406\
        );

    \I__1393\ : Span4Mux_v
    port map (
            O => \N__7436\,
            I => \N__7403\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7433\,
            I => \N__7400\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7428\,
            I => \N__7397\
        );

    \I__1390\ : Span4Mux_h
    port map (
            O => \N__7421\,
            I => \N__7390\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__7418\,
            I => \N__7390\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7415\,
            I => \N__7390\
        );

    \I__1387\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7387\
        );

    \I__1386\ : Sp12to4
    port map (
            O => \N__7411\,
            I => \N__7382\
        );

    \I__1385\ : Sp12to4
    port map (
            O => \N__7406\,
            I => \N__7382\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__7403\,
            I => \N__7379\
        );

    \I__1383\ : Span4Mux_v
    port map (
            O => \N__7400\,
            I => \N__7370\
        );

    \I__1382\ : Span4Mux_h
    port map (
            O => \N__7397\,
            I => \N__7370\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__7390\,
            I => \N__7370\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7370\
        );

    \I__1379\ : Span12Mux_h
    port map (
            O => \N__7382\,
            I => \N__7367\
        );

    \I__1378\ : Span4Mux_v
    port map (
            O => \N__7379\,
            I => \N__7364\
        );

    \I__1377\ : Sp12to4
    port map (
            O => \N__7370\,
            I => \N__7361\
        );

    \I__1376\ : Span12Mux_v
    port map (
            O => \N__7367\,
            I => \N__7358\
        );

    \I__1375\ : Sp12to4
    port map (
            O => \N__7364\,
            I => \N__7353\
        );

    \I__1374\ : Span12Mux_v
    port map (
            O => \N__7361\,
            I => \N__7353\
        );

    \I__1373\ : Odrv12
    port map (
            O => \N__7358\,
            I => \A_c_22\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__7353\,
            I => \A_c_22\
        );

    \I__1371\ : CascadeMux
    port map (
            O => \N__7348\,
            I => \N__7345\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7345\,
            I => \N__7339\
        );

    \I__1369\ : InMux
    port map (
            O => \N__7344\,
            I => \N__7336\
        );

    \I__1368\ : InMux
    port map (
            O => \N__7343\,
            I => \N__7331\
        );

    \I__1367\ : InMux
    port map (
            O => \N__7342\,
            I => \N__7331\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7339\,
            I => \ATA_BASE_0\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__7336\,
            I => \ATA_BASE_0\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7331\,
            I => \ATA_BASE_0\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7324\,
            I => \N__7319\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7323\,
            I => \N__7315\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7322\,
            I => \N__7312\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7309\
        );

    \I__1359\ : InMux
    port map (
            O => \N__7318\,
            I => \N__7306\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__7315\,
            I => \ATA_BASE_6\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7312\,
            I => \ATA_BASE_6\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7309\,
            I => \ATA_BASE_6\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7306\,
            I => \ATA_BASE_6\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7279\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7279\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7279\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7279\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7279\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7292\,
            I => \N__7279\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7279\,
            I => \N__7274\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7278\,
            I => \N__7271\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__7277\,
            I => \N__7268\
        );

    \I__1345\ : Span4Mux_v
    port map (
            O => \N__7274\,
            I => \N__7261\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7271\,
            I => \N__7258\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7247\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7267\,
            I => \N__7247\
        );

    \I__1341\ : InMux
    port map (
            O => \N__7266\,
            I => \N__7247\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7265\,
            I => \N__7247\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7264\,
            I => \N__7247\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__7261\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__7258\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7247\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1335\ : InMux
    port map (
            O => \N__7240\,
            I => \N__7237\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7237\,
            I => \N__7231\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7236\,
            I => \N__7224\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7235\,
            I => \N__7224\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7234\,
            I => \N__7224\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__7231\,
            I => \U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__7224\,
            I => \U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__7219\,
            I => \N__7214\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7209\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7217\,
            I => \N__7209\
        );

    \I__1325\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7206\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7209\,
            I => \N__7203\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7200\
        );

    \I__1322\ : Span4Mux_v
    port map (
            O => \N__7203\,
            I => \N__7195\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__7200\,
            I => \N__7195\
        );

    \I__1320\ : Sp12to4
    port map (
            O => \N__7195\,
            I => \N__7192\
        );

    \I__1319\ : Span12Mux_h
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1318\ : Odrv12
    port map (
            O => \N__7189\,
            I => \D_in_7\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__7186\,
            I => \N__7181\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7178\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7184\,
            I => \N__7175\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7172\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7178\,
            I => \ATA_BASE_3\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7175\,
            I => \ATA_BASE_3\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7172\,
            I => \ATA_BASE_3\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__7165\,
            I => \N__7162\
        );

    \I__1309\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7159\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__7159\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_d\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7153\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__7153\,
            I => \N__7150\
        );

    \I__1305\ : Odrv4
    port map (
            O => \N__7150\,
            I => \U409_ADDRESS_DECODE.g0_i_0Z0Z_0\
        );

    \I__1304\ : InMux
    port map (
            O => \N__7147\,
            I => \N__7144\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__7141\,
            I => \U409_ADDRESS_DECODE.g0_i_o4Z0Z_1\
        );

    \I__1301\ : InMux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__7135\,
            I => \U409_ADDRESS_DECODE.g0_i_o4Z0Z_0\
        );

    \I__1299\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7129\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7129\,
            I => \U409_ADDRESS_DECODE_ATA_ROM_0_1\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__7126\,
            I => \N__7122\
        );

    \I__1296\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7117\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7122\,
            I => \N__7117\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__7117\,
            I => \N__7114\
        );

    \I__1293\ : Odrv4
    port map (
            O => \N__7114\,
            I => \U409_TRANSFER_ACK.CO1\
        );

    \I__1292\ : InMux
    port map (
            O => \N__7111\,
            I => \N__7106\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7103\
        );

    \I__1290\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7100\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7106\,
            I => \N__7096\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7093\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__7100\,
            I => \N__7090\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7087\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__7096\,
            I => \N__7076\
        );

    \I__1284\ : Span4Mux_v
    port map (
            O => \N__7093\,
            I => \N__7076\
        );

    \I__1283\ : Span4Mux_v
    port map (
            O => \N__7090\,
            I => \N__7076\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7087\,
            I => \N__7076\
        );

    \I__1281\ : InMux
    port map (
            O => \N__7086\,
            I => \N__7073\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__7085\,
            I => \N__7070\
        );

    \I__1279\ : Span4Mux_v
    port map (
            O => \N__7076\,
            I => \N__7065\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__7073\,
            I => \N__7065\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7062\
        );

    \I__1276\ : Span4Mux_v
    port map (
            O => \N__7065\,
            I => \N__7059\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__7062\,
            I => \N__7056\
        );

    \I__1274\ : Span4Mux_v
    port map (
            O => \N__7059\,
            I => \N__7053\
        );

    \I__1273\ : Span12Mux_h
    port map (
            O => \N__7056\,
            I => \N__7050\
        );

    \I__1272\ : IoSpan4Mux
    port map (
            O => \N__7053\,
            I => \N__7047\
        );

    \I__1271\ : Odrv12
    port map (
            O => \N__7050\,
            I => \TM_c_1\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__7047\,
            I => \TM_c_1\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__7042\,
            I => \N__7037\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7041\,
            I => \N__7034\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7040\,
            I => \N__7031\
        );

    \I__1266\ : InMux
    port map (
            O => \N__7037\,
            I => \N__7026\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7034\,
            I => \N__7023\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7031\,
            I => \N__7020\
        );

    \I__1263\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7017\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7014\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__7026\,
            I => \N__7010\
        );

    \I__1260\ : Span4Mux_v
    port map (
            O => \N__7023\,
            I => \N__7001\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__7020\,
            I => \N__7001\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__7017\,
            I => \N__7001\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__7014\,
            I => \N__7001\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7013\,
            I => \N__6998\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__7010\,
            I => \N__6995\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__7001\,
            I => \N__6990\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6990\
        );

    \I__1252\ : Sp12to4
    port map (
            O => \N__6995\,
            I => \N__6987\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__6990\,
            I => \N__6984\
        );

    \I__1250\ : Span12Mux_h
    port map (
            O => \N__6987\,
            I => \N__6981\
        );

    \I__1249\ : Span4Mux_v
    port map (
            O => \N__6984\,
            I => \N__6978\
        );

    \I__1248\ : Span12Mux_v
    port map (
            O => \N__6981\,
            I => \N__6975\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__6978\,
            I => \N__6972\
        );

    \I__1246\ : Odrv12
    port map (
            O => \N__6975\,
            I => \TM_c_0\
        );

    \I__1245\ : Odrv4
    port map (
            O => \N__6972\,
            I => \TM_c_0\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6961\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__1241\ : Odrv12
    port map (
            O => \N__6958\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6952\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6952\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__6949\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6946\,
            I => \N__6941\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6945\,
            I => \N__6936\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6936\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6941\,
            I => \ATA_BASE_2\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6936\,
            I => \ATA_BASE_2\
        );

    \I__1232\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \N__6927\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__6930\,
            I => \N__6923\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6920\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6915\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6915\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6912\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6915\,
            I => \N__6909\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__6912\,
            I => \N__6906\
        );

    \I__1224\ : Span4Mux_v
    port map (
            O => \N__6909\,
            I => \N__6903\
        );

    \I__1223\ : Sp12to4
    port map (
            O => \N__6906\,
            I => \N__6900\
        );

    \I__1222\ : Sp12to4
    port map (
            O => \N__6903\,
            I => \N__6895\
        );

    \I__1221\ : Span12Mux_h
    port map (
            O => \N__6900\,
            I => \N__6895\
        );

    \I__1220\ : Odrv12
    port map (
            O => \N__6895\,
            I => \D_in_4\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6888\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \N__6885\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6880\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6880\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6880\,
            I => \N__6877\
        );

    \I__1214\ : Span4Mux_h
    port map (
            O => \N__6877\,
            I => \N__6874\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__6874\,
            I => \N__6870\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6867\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__6870\,
            I => \N__6864\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6867\,
            I => \N__6861\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__6864\,
            I => \N__6858\
        );

    \I__1208\ : Span12Mux_v
    port map (
            O => \N__6861\,
            I => \N__6855\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__6858\,
            I => \D_in_5\
        );

    \I__1206\ : Odrv12
    port map (
            O => \N__6855\,
            I => \D_in_5\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6847\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6847\,
            I => \N__6843\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__6846\,
            I => \N__6840\
        );

    \I__1202\ : Span4Mux_v
    port map (
            O => \N__6843\,
            I => \N__6837\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6833\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__6837\,
            I => \N__6830\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6827\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6833\,
            I => \N__6824\
        );

    \I__1197\ : Sp12to4
    port map (
            O => \N__6830\,
            I => \N__6821\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6818\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6824\,
            I => \N__6815\
        );

    \I__1194\ : Span12Mux_h
    port map (
            O => \N__6821\,
            I => \N__6808\
        );

    \I__1193\ : Span12Mux_v
    port map (
            O => \N__6818\,
            I => \N__6808\
        );

    \I__1192\ : Sp12to4
    port map (
            O => \N__6815\,
            I => \N__6808\
        );

    \I__1191\ : Odrv12
    port map (
            O => \N__6808\,
            I => \D_in_6\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6805\,
            I => \N__6797\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6804\,
            I => \N__6797\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6803\,
            I => \N__6792\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6802\,
            I => \N__6792\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__6797\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6792\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6787\,
            I => \N__6783\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__6786\,
            I => \N__6779\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6783\,
            I => \N__6773\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6770\
        );

    \I__1180\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6765\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6765\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6760\
        );

    \I__1177\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6760\
        );

    \I__1176\ : Span4Mux_h
    port map (
            O => \N__6773\,
            I => \N__6757\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__6770\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6765\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__6760\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__6757\,
            I => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6744\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__6747\,
            I => \N__6741\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__6744\,
            I => \N__6738\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6735\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__6738\,
            I => \BRIDGE_BASE_3\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6735\,
            I => \BRIDGE_BASE_3\
        );

    \I__1165\ : IoInMux
    port map (
            O => \N__6730\,
            I => \N__6727\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6727\,
            I => \N__6724\
        );

    \I__1163\ : Span4Mux_s1_v
    port map (
            O => \N__6724\,
            I => \N__6721\
        );

    \I__1162\ : Sp12to4
    port map (
            O => \N__6721\,
            I => \N__6718\
        );

    \I__1161\ : Span12Mux_h
    port map (
            O => \N__6718\,
            I => \N__6711\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6717\,
            I => \N__6707\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6716\,
            I => \N__6704\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6715\,
            I => \N__6699\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6714\,
            I => \N__6699\
        );

    \I__1156\ : Span12Mux_v
    port map (
            O => \N__6711\,
            I => \N__6695\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6692\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6707\,
            I => \N__6687\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6704\,
            I => \N__6687\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6699\,
            I => \N__6684\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6698\,
            I => \N__6681\
        );

    \I__1150\ : Odrv12
    port map (
            O => \N__6695\,
            I => \CONFIGENn_c\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__6692\,
            I => \CONFIGENn_c\
        );

    \I__1148\ : Odrv12
    port map (
            O => \N__6687\,
            I => \CONFIGENn_c\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__6684\,
            I => \CONFIGENn_c\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6681\,
            I => \CONFIGENn_c\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__6670\,
            I => \N__6666\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6663\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6660\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6663\,
            I => \N__6653\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6653\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6650\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6647\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__6653\,
            I => \ATA_BASE_5\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6650\,
            I => \ATA_BASE_5\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6647\,
            I => \ATA_BASE_5\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6637\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6631\,
            I => \N__6628\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__6628\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6622\,
            I => \N__6616\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6611\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6611\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6608\
        );

    \I__1125\ : Span4Mux_h
    port map (
            O => \N__6616\,
            I => \N__6604\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6611\,
            I => \N__6599\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6608\,
            I => \N__6599\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6607\,
            I => \N__6596\
        );

    \I__1121\ : Span4Mux_v
    port map (
            O => \N__6604\,
            I => \N__6589\
        );

    \I__1120\ : Span4Mux_h
    port map (
            O => \N__6599\,
            I => \N__6589\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6596\,
            I => \N__6589\
        );

    \I__1118\ : Span4Mux_h
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__6583\,
            I => \A_c_31\
        );

    \I__1115\ : IoInMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1113\ : Span12Mux_s9_h
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1112\ : Span12Mux_h
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__6568\,
            I => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6565\,
            I => \N__6561\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6564\,
            I => \N__6558\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6561\,
            I => \N__6555\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6552\
        );

    \I__1106\ : Span4Mux_v
    port map (
            O => \N__6555\,
            I => \N__6549\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__6552\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__6549\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__6544\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6538\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__6538\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\
        );

    \I__1100\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6532\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6532\,
            I => \U409_ADDRESS_DECODE.g2Z0Z_5\
        );

    \I__1098\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6524\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6521\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6518\
        );

    \I__1095\ : LocalMux
    port map (
            O => \N__6524\,
            I => \N__6514\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6521\,
            I => \N__6511\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6518\,
            I => \N__6508\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6517\,
            I => \N__6504\
        );

    \I__1091\ : Span4Mux_h
    port map (
            O => \N__6514\,
            I => \N__6499\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__6511\,
            I => \N__6499\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__6508\,
            I => \N__6496\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6507\,
            I => \N__6493\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6504\,
            I => \N__6490\
        );

    \I__1086\ : Span4Mux_v
    port map (
            O => \N__6499\,
            I => \N__6487\
        );

    \I__1085\ : Span4Mux_v
    port map (
            O => \N__6496\,
            I => \N__6482\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6482\
        );

    \I__1083\ : Sp12to4
    port map (
            O => \N__6490\,
            I => \N__6479\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__6487\,
            I => \N__6476\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__6482\,
            I => \N__6473\
        );

    \I__1080\ : Span12Mux_v
    port map (
            O => \N__6479\,
            I => \N__6470\
        );

    \I__1079\ : Sp12to4
    port map (
            O => \N__6476\,
            I => \N__6465\
        );

    \I__1078\ : Span12Mux_v
    port map (
            O => \N__6473\,
            I => \N__6465\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__6470\,
            I => \A_c_28\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__6465\,
            I => \A_c_28\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U409_ADDRESS_DECODE_g2_6\
        );

    \I__1073\ : CascadeMux
    port map (
            O => \N__6454\,
            I => \U409_ADDRESS_DECODE_g2_7_cascade_\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__6445\,
            I => \U409_TRANSFER_ACK.G_14_0_o7_0\
        );

    \I__1069\ : IoInMux
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__1067\ : Span4Mux_s0_h
    port map (
            O => \N__6436\,
            I => \N__6433\
        );

    \I__1066\ : Sp12to4
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1065\ : Span12Mux_s11_v
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1064\ : Span12Mux_h
    port map (
            O => \N__6427\,
            I => \N__6424\
        );

    \I__1063\ : Odrv12
    port map (
            O => \N__6424\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__6418\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__6412\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__6409\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6397\
        );

    \I__1055\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6391\
        );

    \I__1054\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6391\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6388\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6397\,
            I => \N__6384\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6396\,
            I => \N__6381\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6376\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6388\,
            I => \N__6376\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6387\,
            I => \N__6373\
        );

    \I__1047\ : Span4Mux_v
    port map (
            O => \N__6384\,
            I => \N__6367\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6381\,
            I => \N__6367\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__6376\,
            I => \N__6364\
        );

    \I__1044\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6361\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6358\
        );

    \I__1042\ : Span4Mux_v
    port map (
            O => \N__6367\,
            I => \N__6355\
        );

    \I__1041\ : Sp12to4
    port map (
            O => \N__6364\,
            I => \N__6348\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6348\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6358\,
            I => \N__6348\
        );

    \I__1038\ : Sp12to4
    port map (
            O => \N__6355\,
            I => \N__6345\
        );

    \I__1037\ : Span12Mux_h
    port map (
            O => \N__6348\,
            I => \N__6342\
        );

    \I__1036\ : Span12Mux_h
    port map (
            O => \N__6345\,
            I => \N__6339\
        );

    \I__1035\ : Span12Mux_v
    port map (
            O => \N__6342\,
            I => \N__6336\
        );

    \I__1034\ : Span12Mux_v
    port map (
            O => \N__6339\,
            I => \N__6333\
        );

    \I__1033\ : Odrv12
    port map (
            O => \N__6336\,
            I => \RnW_c\
        );

    \I__1032\ : Odrv12
    port map (
            O => \N__6333\,
            I => \RnW_c\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6328\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1028\ : Odrv4
    port map (
            O => \N__6319\,
            I => \U409_ADDRESS_DECODE.g2Z0Z_10\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \U409_ADDRESS_DECODE.g2Z0Z_11_cascade_\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__6304\,
            I => \U409_ADDRESS_DECODE.g2Z0Z_9\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6289\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6289\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__6299\,
            I => \N__6285\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__6298\,
            I => \N__6282\
        );

    \I__1018\ : CascadeMux
    port map (
            O => \N__6297\,
            I => \N__6279\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__6296\,
            I => \N__6276\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6271\
        );

    \I__1015\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6271\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6267\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6262\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6262\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6257\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6279\,
            I => \N__6257\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6254\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6271\,
            I => \N__6251\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6270\,
            I => \N__6248\
        );

    \I__1006\ : Span4Mux_h
    port map (
            O => \N__6267\,
            I => \N__6234\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6234\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__6257\,
            I => \N__6234\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6234\
        );

    \I__1002\ : Span4Mux_v
    port map (
            O => \N__6251\,
            I => \N__6228\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__6248\,
            I => \N__6228\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6221\
        );

    \I__999\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6221\
        );

    \I__998\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6221\
        );

    \I__997\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6216\
        );

    \I__996\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6216\
        );

    \I__995\ : Span4Mux_v
    port map (
            O => \N__6234\,
            I => \N__6213\
        );

    \I__994\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6210\
        );

    \I__993\ : Span4Mux_h
    port map (
            O => \N__6228\,
            I => \N__6203\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6203\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__6216\,
            I => \N__6203\
        );

    \I__990\ : Sp12to4
    port map (
            O => \N__6213\,
            I => \N__6198\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6210\,
            I => \N__6198\
        );

    \I__988\ : Span4Mux_v
    port map (
            O => \N__6203\,
            I => \N__6195\
        );

    \I__987\ : Span12Mux_h
    port map (
            O => \N__6198\,
            I => \N__6192\
        );

    \I__986\ : Span4Mux_h
    port map (
            O => \N__6195\,
            I => \N__6189\
        );

    \I__985\ : Span12Mux_v
    port map (
            O => \N__6192\,
            I => \N__6186\
        );

    \I__984\ : Sp12to4
    port map (
            O => \N__6189\,
            I => \N__6183\
        );

    \I__983\ : Odrv12
    port map (
            O => \N__6186\,
            I => \A_c_1\
        );

    \I__982\ : Odrv12
    port map (
            O => \N__6183\,
            I => \A_c_1\
        );

    \I__981\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6171\
        );

    \I__980\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6171\
        );

    \I__979\ : InMux
    port map (
            O => \N__6176\,
            I => \N__6167\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6164\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6170\,
            I => \N__6161\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6155\
        );

    \I__975\ : Span4Mux_v
    port map (
            O => \N__6164\,
            I => \N__6151\
        );

    \I__974\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6148\
        );

    \I__973\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6145\
        );

    \I__972\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6140\
        );

    \I__971\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6140\
        );

    \I__970\ : Span4Mux_h
    port map (
            O => \N__6155\,
            I => \N__6137\
        );

    \I__969\ : InMux
    port map (
            O => \N__6154\,
            I => \N__6134\
        );

    \I__968\ : Odrv4
    port map (
            O => \N__6151\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6148\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6145\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6140\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__964\ : Odrv4
    port map (
            O => \N__6137\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6134\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__962\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6115\
        );

    \I__961\ : InMux
    port map (
            O => \N__6120\,
            I => \N__6115\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__6115\,
            I => \N__6112\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__6112\,
            I => \U409_AUTOCONFIG.un1_STATE_1_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6105\
        );

    \I__957\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6102\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6105\,
            I => \N__6099\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6102\,
            I => \N__6096\
        );

    \I__954\ : Odrv4
    port map (
            O => \N__6099\,
            I => \BRIDGE_BASE_0\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__6096\,
            I => \BRIDGE_BASE_0\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__6091\,
            I => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_\
        );

    \I__951\ : InMux
    port map (
            O => \N__6088\,
            I => \N__6082\
        );

    \I__950\ : InMux
    port map (
            O => \N__6087\,
            I => \N__6082\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6082\,
            I => \N__6078\
        );

    \I__948\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6075\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__6078\,
            I => \N__6071\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__6075\,
            I => \N__6068\
        );

    \I__945\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6065\
        );

    \I__944\ : Span4Mux_v
    port map (
            O => \N__6071\,
            I => \N__6062\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__6068\,
            I => \N__6059\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6065\,
            I => \N__6056\
        );

    \I__941\ : Span4Mux_h
    port map (
            O => \N__6062\,
            I => \N__6053\
        );

    \I__940\ : Span4Mux_v
    port map (
            O => \N__6059\,
            I => \N__6050\
        );

    \I__939\ : Sp12to4
    port map (
            O => \N__6056\,
            I => \N__6047\
        );

    \I__938\ : Sp12to4
    port map (
            O => \N__6053\,
            I => \N__6040\
        );

    \I__937\ : Sp12to4
    port map (
            O => \N__6050\,
            I => \N__6040\
        );

    \I__936\ : Span12Mux_v
    port map (
            O => \N__6047\,
            I => \N__6040\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__6040\,
            I => \A_c_26\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \N__6033\
        );

    \I__933\ : InMux
    port map (
            O => \N__6036\,
            I => \N__6027\
        );

    \I__932\ : InMux
    port map (
            O => \N__6033\,
            I => \N__6027\
        );

    \I__931\ : InMux
    port map (
            O => \N__6032\,
            I => \N__6023\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6027\,
            I => \N__6020\
        );

    \I__929\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6017\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__6014\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__6020\,
            I => \N__6011\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__6008\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__6014\,
            I => \N__6005\
        );

    \I__924\ : Span4Mux_h
    port map (
            O => \N__6011\,
            I => \N__6000\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__6008\,
            I => \N__6000\
        );

    \I__922\ : Sp12to4
    port map (
            O => \N__6005\,
            I => \N__5995\
        );

    \I__921\ : Sp12to4
    port map (
            O => \N__6000\,
            I => \N__5995\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__5995\,
            I => \A_c_25\
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__5992\,
            I => \N__5988\
        );

    \I__918\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5984\
        );

    \I__917\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5979\
        );

    \I__916\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5979\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5984\,
            I => \N__5975\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5979\,
            I => \N__5972\
        );

    \I__913\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5969\
        );

    \I__912\ : Span4Mux_v
    port map (
            O => \N__5975\,
            I => \N__5966\
        );

    \I__911\ : Span4Mux_h
    port map (
            O => \N__5972\,
            I => \N__5963\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__5969\,
            I => \N__5960\
        );

    \I__909\ : Span4Mux_v
    port map (
            O => \N__5966\,
            I => \N__5957\
        );

    \I__908\ : Sp12to4
    port map (
            O => \N__5963\,
            I => \N__5952\
        );

    \I__907\ : Sp12to4
    port map (
            O => \N__5960\,
            I => \N__5952\
        );

    \I__906\ : Sp12to4
    port map (
            O => \N__5957\,
            I => \N__5947\
        );

    \I__905\ : Span12Mux_v
    port map (
            O => \N__5952\,
            I => \N__5947\
        );

    \I__904\ : Odrv12
    port map (
            O => \N__5947\,
            I => \A_c_24\
        );

    \I__903\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5941\,
            I => \U409_ADDRESS_DECODE.g2Z0Z_4\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__5938\,
            I => \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_\
        );

    \I__900\ : CascadeMux
    port map (
            O => \N__5935\,
            I => \N__5931\
        );

    \I__899\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5928\
        );

    \I__898\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5925\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__5928\,
            I => \N__5917\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5925\,
            I => \N__5917\
        );

    \I__895\ : InMux
    port map (
            O => \N__5924\,
            I => \N__5914\
        );

    \I__894\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5911\
        );

    \I__893\ : InMux
    port map (
            O => \N__5922\,
            I => \N__5908\
        );

    \I__892\ : Odrv4
    port map (
            O => \N__5917\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__5914\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5911\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5908\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__888\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5895\
        );

    \I__887\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5892\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__5895\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5892\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__884\ : CascadeMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__883\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5880\
        );

    \I__882\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5877\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5880\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__5877\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__879\ : IoInMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__877\ : IoSpan4Mux
    port map (
            O => \N__5866\,
            I => \N__5863\
        );

    \I__876\ : Span4Mux_s2_v
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__875\ : Sp12to4
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__874\ : Span12Mux_s11_v
    port map (
            O => \N__5857\,
            I => \N__5854\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__5854\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_2\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__5851\,
            I => \N__5848\
        );

    \I__871\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5845\,
            I => \N__5841\
        );

    \I__869\ : InMux
    port map (
            O => \N__5844\,
            I => \N__5838\
        );

    \I__868\ : Odrv12
    port map (
            O => \N__5841\,
            I => \BRIDGE_BASE_1\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5838\,
            I => \BRIDGE_BASE_1\
        );

    \I__866\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__5830\,
            I => \N__5826\
        );

    \I__864\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5823\
        );

    \I__863\ : Odrv12
    port map (
            O => \N__5826\,
            I => \BRIDGE_BASE_2\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5823\,
            I => \BRIDGE_BASE_2\
        );

    \I__861\ : InMux
    port map (
            O => \N__5818\,
            I => \N__5811\
        );

    \I__860\ : InMux
    port map (
            O => \N__5817\,
            I => \N__5803\
        );

    \I__859\ : InMux
    port map (
            O => \N__5816\,
            I => \N__5803\
        );

    \I__858\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5803\
        );

    \I__857\ : InMux
    port map (
            O => \N__5814\,
            I => \N__5799\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5796\
        );

    \I__855\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5793\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5790\
        );

    \I__853\ : CascadeMux
    port map (
            O => \N__5802\,
            I => \N__5785\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__5799\,
            I => \N__5782\
        );

    \I__851\ : Sp12to4
    port map (
            O => \N__5796\,
            I => \N__5777\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5793\,
            I => \N__5777\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__5790\,
            I => \N__5774\
        );

    \I__848\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5771\
        );

    \I__847\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5768\
        );

    \I__846\ : InMux
    port map (
            O => \N__5785\,
            I => \N__5765\
        );

    \I__845\ : Span12Mux_v
    port map (
            O => \N__5782\,
            I => \N__5762\
        );

    \I__844\ : Span12Mux_v
    port map (
            O => \N__5777\,
            I => \N__5751\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__5774\,
            I => \N__5751\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__5771\,
            I => \N__5751\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5768\,
            I => \N__5751\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__5765\,
            I => \N__5751\
        );

    \I__839\ : Odrv12
    port map (
            O => \N__5762\,
            I => \A_c_5\
        );

    \I__838\ : Odrv12
    port map (
            O => \N__5751\,
            I => \A_c_5\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5746\,
            I => \N__5742\
        );

    \I__836\ : InMux
    port map (
            O => \N__5745\,
            I => \N__5737\
        );

    \I__835\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5737\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U409_AUTOCONFIG.N_68\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__5734\,
            I => \N__5730\
        );

    \I__832\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5724\
        );

    \I__831\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5721\
        );

    \I__830\ : InMux
    port map (
            O => \N__5729\,
            I => \N__5716\
        );

    \I__829\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5716\
        );

    \I__828\ : InMux
    port map (
            O => \N__5727\,
            I => \N__5713\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__5724\,
            I => \N__5709\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5704\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5704\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__5713\,
            I => \N__5698\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__5712\,
            I => \N__5690\
        );

    \I__822\ : Span4Mux_v
    port map (
            O => \N__5709\,
            I => \N__5685\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__5704\,
            I => \N__5685\
        );

    \I__820\ : InMux
    port map (
            O => \N__5703\,
            I => \N__5680\
        );

    \I__819\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5680\
        );

    \I__818\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5677\
        );

    \I__817\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5674\
        );

    \I__816\ : InMux
    port map (
            O => \N__5697\,
            I => \N__5667\
        );

    \I__815\ : InMux
    port map (
            O => \N__5696\,
            I => \N__5667\
        );

    \I__814\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5667\
        );

    \I__813\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5664\
        );

    \I__812\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5659\
        );

    \I__811\ : InMux
    port map (
            O => \N__5690\,
            I => \N__5659\
        );

    \I__810\ : Sp12to4
    port map (
            O => \N__5685\,
            I => \N__5644\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5644\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5644\
        );

    \I__807\ : Sp12to4
    port map (
            O => \N__5674\,
            I => \N__5644\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5667\,
            I => \N__5644\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5664\,
            I => \N__5644\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5644\
        );

    \I__803\ : Odrv12
    port map (
            O => \N__5644\,
            I => \A_c_4\
        );

    \I__802\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5638\,
            I => \U409_AUTOCONFIG.N_47\
        );

    \I__800\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__797\ : Sp12to4
    port map (
            O => \N__5626\,
            I => \N__5623\
        );

    \I__796\ : Span12Mux_h
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__795\ : Span12Mux_h
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__794\ : Span12Mux_v
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__5614\,
            I => \AUTOBOOT_c\
        );

    \I__792\ : InMux
    port map (
            O => \N__5611\,
            I => \N__5607\
        );

    \I__791\ : InMux
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5607\,
            I => \N__5601\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5604\,
            I => \N__5598\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__5601\,
            I => \N__5594\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__5598\,
            I => \N__5591\
        );

    \I__786\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5588\
        );

    \I__785\ : Odrv4
    port map (
            O => \N__5594\,
            I => \U409_AUTOCONFIG.N_196_1\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__5591\,
            I => \U409_AUTOCONFIG.N_196_1\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__5588\,
            I => \U409_AUTOCONFIG.N_196_1\
        );

    \I__782\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5570\
        );

    \I__781\ : InMux
    port map (
            O => \N__5580\,
            I => \N__5570\
        );

    \I__780\ : InMux
    port map (
            O => \N__5579\,
            I => \N__5565\
        );

    \I__779\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5565\
        );

    \I__778\ : InMux
    port map (
            O => \N__5577\,
            I => \N__5561\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__5576\,
            I => \N__5556\
        );

    \I__776\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5552\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5570\,
            I => \N__5547\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5565\,
            I => \N__5547\
        );

    \I__773\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5544\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__5561\,
            I => \N__5537\
        );

    \I__771\ : InMux
    port map (
            O => \N__5560\,
            I => \N__5534\
        );

    \I__770\ : InMux
    port map (
            O => \N__5559\,
            I => \N__5531\
        );

    \I__769\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5526\
        );

    \I__768\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5526\
        );

    \I__767\ : InMux
    port map (
            O => \N__5552\,
            I => \N__5523\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__5547\,
            I => \N__5518\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5518\
        );

    \I__764\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5513\
        );

    \I__763\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5513\
        );

    \I__762\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5508\
        );

    \I__761\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5508\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__5537\,
            I => \N__5501\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5501\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5501\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__5526\,
            I => \N__5498\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5523\,
            I => \N__5495\
        );

    \I__755\ : Span4Mux_h
    port map (
            O => \N__5518\,
            I => \N__5488\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5488\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5508\,
            I => \N__5488\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__5501\,
            I => \N__5485\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__5498\,
            I => \N__5478\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__5495\,
            I => \N__5478\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__5488\,
            I => \N__5478\
        );

    \I__748\ : Sp12to4
    port map (
            O => \N__5485\,
            I => \N__5473\
        );

    \I__747\ : Sp12to4
    port map (
            O => \N__5478\,
            I => \N__5473\
        );

    \I__746\ : Span12Mux_h
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__5470\,
            I => \A_c_2\
        );

    \I__744\ : InMux
    port map (
            O => \N__5467\,
            I => \N__5459\
        );

    \I__743\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5459\
        );

    \I__742\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5456\
        );

    \I__741\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \N__5452\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5459\,
            I => \N__5445\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5456\,
            I => \N__5442\
        );

    \I__738\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5437\
        );

    \I__737\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5437\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__5451\,
            I => \N__5434\
        );

    \I__735\ : InMux
    port map (
            O => \N__5450\,
            I => \N__5428\
        );

    \I__734\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5425\
        );

    \I__733\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5422\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__5445\,
            I => \N__5419\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__5442\,
            I => \N__5414\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5437\,
            I => \N__5414\
        );

    \I__729\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5409\
        );

    \I__728\ : InMux
    port map (
            O => \N__5433\,
            I => \N__5409\
        );

    \I__727\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5406\
        );

    \I__726\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5403\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__5428\,
            I => \N__5400\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5425\,
            I => \N__5387\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5422\,
            I => \N__5387\
        );

    \I__722\ : Sp12to4
    port map (
            O => \N__5419\,
            I => \N__5387\
        );

    \I__721\ : Sp12to4
    port map (
            O => \N__5414\,
            I => \N__5387\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5409\,
            I => \N__5387\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5406\,
            I => \N__5387\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5384\
        );

    \I__717\ : Sp12to4
    port map (
            O => \N__5400\,
            I => \N__5381\
        );

    \I__716\ : Span12Mux_h
    port map (
            O => \N__5387\,
            I => \N__5378\
        );

    \I__715\ : Span12Mux_v
    port map (
            O => \N__5384\,
            I => \N__5375\
        );

    \I__714\ : Span12Mux_v
    port map (
            O => \N__5381\,
            I => \N__5372\
        );

    \I__713\ : Span12Mux_v
    port map (
            O => \N__5378\,
            I => \N__5369\
        );

    \I__712\ : Odrv12
    port map (
            O => \N__5375\,
            I => \A_c_3\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__5372\,
            I => \A_c_3\
        );

    \I__710\ : Odrv12
    port map (
            O => \N__5369\,
            I => \A_c_3\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__708\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5356\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5356\,
            I => \N__5353\
        );

    \I__706\ : Odrv4
    port map (
            O => \N__5353\,
            I => \U409_AUTOCONFIG.N_54\
        );

    \I__705\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5347\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5347\,
            I => \U409_ADDRESS_DECODE.g2_5_0\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__5344\,
            I => \U409_ADDRESS_DECODE.g2_6_0_cascade_\
        );

    \I__702\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__701\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5329\
        );

    \I__700\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5329\
        );

    \I__699\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5326\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5335\,
            I => \N__5323\
        );

    \I__697\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5320\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5329\,
            I => \N__5315\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5315\
        );

    \I__694\ : Span4Mux_v
    port map (
            O => \N__5323\,
            I => \N__5312\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5307\
        );

    \I__692\ : Sp12to4
    port map (
            O => \N__5315\,
            I => \N__5307\
        );

    \I__691\ : Span4Mux_v
    port map (
            O => \N__5312\,
            I => \N__5304\
        );

    \I__690\ : Span12Mux_v
    port map (
            O => \N__5307\,
            I => \N__5301\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__5304\,
            I => \N__5298\
        );

    \I__688\ : Odrv12
    port map (
            O => \N__5301\,
            I => \A_c_29\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__5298\,
            I => \A_c_29\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__5293\,
            I => \N__5288\
        );

    \I__685\ : InMux
    port map (
            O => \N__5292\,
            I => \N__5283\
        );

    \I__684\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5283\
        );

    \I__683\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5280\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5283\,
            I => \N__5275\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5272\
        );

    \I__680\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5269\
        );

    \I__679\ : InMux
    port map (
            O => \N__5278\,
            I => \N__5266\
        );

    \I__678\ : Span4Mux_h
    port map (
            O => \N__5275\,
            I => \N__5259\
        );

    \I__677\ : Span4Mux_h
    port map (
            O => \N__5272\,
            I => \N__5259\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5259\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5266\,
            I => \N__5256\
        );

    \I__674\ : Span4Mux_h
    port map (
            O => \N__5259\,
            I => \N__5253\
        );

    \I__673\ : Span12Mux_v
    port map (
            O => \N__5256\,
            I => \N__5250\
        );

    \I__672\ : Span4Mux_v
    port map (
            O => \N__5253\,
            I => \N__5247\
        );

    \I__671\ : Odrv12
    port map (
            O => \N__5250\,
            I => \A_c_30\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__5247\,
            I => \A_c_30\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__5242\,
            I => \N__5236\
        );

    \I__668\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5231\
        );

    \I__667\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5231\
        );

    \I__666\ : InMux
    port map (
            O => \N__5239\,
            I => \N__5228\
        );

    \I__665\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5225\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5222\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__5228\,
            I => \N__5219\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5216\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__5222\,
            I => \N__5213\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__5219\,
            I => \N__5210\
        );

    \I__659\ : Span4Mux_v
    port map (
            O => \N__5216\,
            I => \N__5207\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__5213\,
            I => \N__5202\
        );

    \I__657\ : Sp12to4
    port map (
            O => \N__5210\,
            I => \N__5202\
        );

    \I__656\ : Sp12to4
    port map (
            O => \N__5207\,
            I => \N__5199\
        );

    \I__655\ : Odrv12
    port map (
            O => \N__5202\,
            I => \A_c_27\
        );

    \I__654\ : Odrv12
    port map (
            O => \N__5199\,
            I => \A_c_27\
        );

    \I__653\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5191\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5191\,
            I => \U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3\
        );

    \I__651\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5185\,
            I => \U409_ADDRESS_DECODE.g0_i_a4Z0Z_1\
        );

    \I__649\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5178\
        );

    \I__648\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5175\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__5178\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__645\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__643\ : Span4Mux_h
    port map (
            O => \N__5164\,
            I => \N__5161\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__5161\,
            I => \U409_AUTOCONFIG.LIDE_OUTc_0_0\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__5158\,
            I => \N__5155\
        );

    \I__640\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5152\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__5152\,
            I => \N__5148\
        );

    \I__638\ : InMux
    port map (
            O => \N__5151\,
            I => \N__5145\
        );

    \I__637\ : Odrv12
    port map (
            O => \N__5148\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5145\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\
        );

    \I__635\ : InMux
    port map (
            O => \N__5140\,
            I => \N__5137\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__5137\,
            I => \U409_AUTOCONFIG.N_50\
        );

    \I__633\ : CascadeMux
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__632\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__5125\,
            I => \U409_AUTOCONFIG.LIDE_OUTc_0_0_0\
        );

    \I__629\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__5119\,
            I => \N__5116\
        );

    \I__627\ : Span4Mux_v
    port map (
            O => \N__5116\,
            I => \N__5112\
        );

    \I__626\ : InMux
    port map (
            O => \N__5115\,
            I => \N__5109\
        );

    \I__625\ : Odrv4
    port map (
            O => \N__5112\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__5109\,
            I => \U409_AUTOCONFIG.N_48\
        );

    \I__623\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5092\
        );

    \I__622\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5092\
        );

    \I__621\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5092\
        );

    \I__620\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5092\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5092\,
            I => \U409_AUTOCONFIG.AC_START_RNI777KZ0Z2\
        );

    \I__618\ : InMux
    port map (
            O => \N__5089\,
            I => \N__5085\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__5088\,
            I => \N__5082\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5079\
        );

    \I__615\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5076\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__5079\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5076\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__612\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5065\
        );

    \I__611\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5065\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__5065\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__609\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5058\
        );

    \I__608\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5055\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5058\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__5055\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1\
        );

    \I__605\ : IoInMux
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__603\ : Span12Mux_s4_v
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__602\ : Span12Mux_v
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__601\ : Odrv12
    port map (
            O => \N__5038\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_1\
        );

    \I__600\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__5028\
        );

    \I__598\ : InMux
    port map (
            O => \N__5031\,
            I => \N__5025\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__5028\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__5025\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__595\ : IoInMux
    port map (
            O => \N__5020\,
            I => \N__5017\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__593\ : Span4Mux_s3_v
    port map (
            O => \N__5014\,
            I => \N__5011\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__5011\,
            I => \N__5008\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__590\ : Odrv4
    port map (
            O => \N__5005\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_0\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__5002\,
            I => \U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_\
        );

    \I__588\ : InMux
    port map (
            O => \N__4999\,
            I => \N__4994\
        );

    \I__587\ : InMux
    port map (
            O => \N__4998\,
            I => \N__4991\
        );

    \I__586\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4988\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4994\,
            I => \N__4981\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4981\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4981\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4981\,
            I => \N__4978\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__4978\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_18\
        );

    \I__580\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4968\
        );

    \I__579\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4968\
        );

    \I__578\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4962\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4959\
        );

    \I__576\ : InMux
    port map (
            O => \N__4967\,
            I => \N__4956\
        );

    \I__575\ : InMux
    port map (
            O => \N__4966\,
            I => \N__4953\
        );

    \I__574\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4950\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4962\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__4959\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4956\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4953\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__4950\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__568\ : CascadeMux
    port map (
            O => \N__4939\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\
        );

    \I__567\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__565\ : Odrv4
    port map (
            O => \N__4930\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4\
        );

    \I__564\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4924\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__4921\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_\
        );

    \I__561\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4915\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__558\ : Span4Mux_v
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__557\ : IoSpan4Mux
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__4903\,
            I => \TT_c_1\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__554\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__552\ : Span4Mux_h
    port map (
            O => \N__4891\,
            I => \N__4888\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__4888\,
            I => \N__4885\
        );

    \I__550\ : Span4Mux_v
    port map (
            O => \N__4885\,
            I => \N__4882\
        );

    \I__549\ : Odrv4
    port map (
            O => \N__4882\,
            I => \TT_c_0\
        );

    \I__548\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4876\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\
        );

    \I__546\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4870\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__4867\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__4864\,
            I => \AUTOCONFIG_SPACE_cascade_\
        );

    \I__542\ : IoInMux
    port map (
            O => \N__4861\,
            I => \N__4858\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__4858\,
            I => \N__4853\
        );

    \I__540\ : IoInMux
    port map (
            O => \N__4857\,
            I => \N__4850\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__4856\,
            I => \N__4847\
        );

    \I__538\ : IoSpan4Mux
    port map (
            O => \N__4853\,
            I => \N__4839\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4839\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4839\
        );

    \I__535\ : IoInMux
    port map (
            O => \N__4846\,
            I => \N__4836\
        );

    \I__534\ : IoSpan4Mux
    port map (
            O => \N__4839\,
            I => \N__4831\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__4836\,
            I => \N__4831\
        );

    \I__532\ : Span4Mux_s3_v
    port map (
            O => \N__4831\,
            I => \N__4828\
        );

    \I__531\ : Span4Mux_v
    port map (
            O => \N__4828\,
            I => \N__4825\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__529\ : Odrv4
    port map (
            O => \N__4822\,
            I => \D_1_i\
        );

    \I__528\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4816\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__4816\,
            I => \N__4813\
        );

    \I__526\ : Odrv12
    port map (
            O => \N__4813\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \N__4807\
        );

    \I__524\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4804\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4804\,
            I => \N__4801\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__4801\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0\
        );

    \I__521\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4791\
        );

    \I__520\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4791\
        );

    \I__519\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4788\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__4791\,
            I => \U409_AUTOCONFIG.N_59_1\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__4788\,
            I => \U409_AUTOCONFIG.N_59_1\
        );

    \I__516\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4780\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__4780\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa\
        );

    \I__514\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__4771\,
            I => \N__4767\
        );

    \I__511\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4764\
        );

    \I__510\ : Sp12to4
    port map (
            O => \N__4767\,
            I => \N__4759\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4759\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__4759\,
            I => \U409_AUTOCONFIG.N_57\
        );

    \I__507\ : InMux
    port map (
            O => \N__4756\,
            I => \N__4753\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4753\,
            I => \N__4750\
        );

    \I__505\ : Span4Mux_h
    port map (
            O => \N__4750\,
            I => \N__4747\
        );

    \I__504\ : Odrv4
    port map (
            O => \N__4747\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1\
        );

    \I__503\ : CascadeMux
    port map (
            O => \N__4744\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__4741\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_\
        );

    \I__501\ : CascadeMux
    port map (
            O => \N__4738\,
            I => \U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__4735\,
            I => \U409_AUTOCONFIG.N_55_cascade_\
        );

    \I__499\ : InMux
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4725\
        );

    \I__497\ : InMux
    port map (
            O => \N__4728\,
            I => \N__4722\
        );

    \I__496\ : Odrv4
    port map (
            O => \N__4725\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4722\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__4717\,
            I => \N__4714\
        );

    \I__493\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4710\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__4713\,
            I => \N__4707\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4710\,
            I => \N__4704\
        );

    \I__490\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4701\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__4704\,
            I => \N__4698\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__4701\,
            I => \N__4695\
        );

    \I__487\ : Sp12to4
    port map (
            O => \N__4698\,
            I => \N__4692\
        );

    \I__486\ : Span4Mux_h
    port map (
            O => \N__4695\,
            I => \N__4689\
        );

    \I__485\ : Span12Mux_s10_h
    port map (
            O => \N__4692\,
            I => \N__4684\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4689\,
            I => \N__4684\
        );

    \I__483\ : Span12Mux_v
    port map (
            O => \N__4684\,
            I => \N__4681\
        );

    \I__482\ : Odrv12
    port map (
            O => \N__4681\,
            I => \CPUCONFn_c\
        );

    \I__481\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4675\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4675\,
            I => \N__4672\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__4672\,
            I => \N__4669\
        );

    \I__478\ : Odrv4
    port map (
            O => \N__4669\,
            I => \U409_AUTOCONFIG.N_40\
        );

    \I__477\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \U409_AUTOCONFIG.N_59_1_cascade_\
        );

    \I__476\ : InMux
    port map (
            O => \N__4663\,
            I => \N__4660\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__4660\,
            I => \N__4656\
        );

    \I__474\ : InMux
    port map (
            O => \N__4659\,
            I => \N__4653\
        );

    \I__473\ : Odrv12
    port map (
            O => \N__4656\,
            I => \U409_AUTOCONFIG.N_61\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4653\,
            I => \U409_AUTOCONFIG.N_61\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__4648\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4639\
        );

    \I__469\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4639\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4639\,
            I => \N__4636\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__4636\,
            I => \U409_AUTOCONFIG.N_67\
        );

    \I__466\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__4630\,
            I => \U409_AUTOCONFIG.N_56\
        );

    \I__464\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4624\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4621\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__4618\,
            I => \N__4615\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__459\ : Span4Mux_h
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__458\ : Odrv4
    port map (
            O => \N__4609\,
            I => \U409_AUTOCONFIG.ATA_BASE10Z0Z_2\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4606\,
            I => \U409_AUTOCONFIG.ATA_BASE10_cascade_\
        );

    \I__456\ : IoInMux
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__454\ : Span12Mux_s2_v
    port map (
            O => \N__4597\,
            I => \N__4594\
        );

    \I__453\ : Span12Mux_v
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__4591\,
            I => \U409_AUTOCONFIG_D_OUT_0_i_3\
        );

    \I__451\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4585\,
            I => \N__4580\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4584\,
            I => \N__4577\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__4583\,
            I => \N__4573\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4580\,
            I => \N__4568\
        );

    \I__446\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4559\
        );

    \I__445\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4559\
        );

    \I__444\ : InMux
    port map (
            O => \N__4573\,
            I => \N__4559\
        );

    \I__443\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4559\
        );

    \I__442\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4556\
        );

    \I__441\ : Sp12to4
    port map (
            O => \N__4568\,
            I => \N__4549\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4559\,
            I => \N__4549\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__4556\,
            I => \N__4549\
        );

    \I__438\ : Odrv12
    port map (
            O => \N__4549\,
            I => \A_c_6\
        );

    \I__437\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4534\
        );

    \I__436\ : InMux
    port map (
            O => \N__4545\,
            I => \N__4534\
        );

    \I__435\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4534\
        );

    \I__434\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4534\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4534\,
            I => \N__4529\
        );

    \I__432\ : InMux
    port map (
            O => \N__4533\,
            I => \N__4526\
        );

    \I__431\ : InMux
    port map (
            O => \N__4532\,
            I => \N__4523\
        );

    \I__430\ : Span4Mux_v
    port map (
            O => \N__4529\,
            I => \N__4520\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4515\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4523\,
            I => \N__4515\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__4520\,
            I => \N__4510\
        );

    \I__426\ : Span12Mux_v
    port map (
            O => \N__4515\,
            I => \N__4510\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4510\,
            I => \A_c_7\
        );

    \I__424\ : CascadeMux
    port map (
            O => \N__4507\,
            I => \U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_\
        );

    \I__423\ : CascadeMux
    port map (
            O => \N__4504\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_\
        );

    \I__422\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__4498\,
            I => \U409_AUTOCONFIG.N_63\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__4495\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \U409_AUTOCONFIG.N_196_1_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4486\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4486\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__4483\,
            I => \U409_AUTOCONFIG.N_67_cascade_\
        );

    \I__415\ : CascadeMux
    port map (
            O => \N__4480\,
            I => \N__4476\
        );

    \I__414\ : InMux
    port map (
            O => \N__4479\,
            I => \N__4473\
        );

    \I__413\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4470\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4473\,
            I => \U409_AUTOCONFIG.N_214_1\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4470\,
            I => \U409_AUTOCONFIG.N_214_1\
        );

    \I__410\ : IoInMux
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__408\ : Span4Mux_s2_h
    port map (
            O => \N__4459\,
            I => \N__4456\
        );

    \I__407\ : Sp12to4
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__406\ : Span12Mux_v
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__405\ : Span12Mux_v
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__404\ : Odrv12
    port map (
            O => \N__4447\,
            I => \PIO_P0_c\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__400\ : Span4Mux_s2_h
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__399\ : Sp12to4
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__398\ : Span12Mux_v
    port map (
            O => \N__4429\,
            I => \N__4426\
        );

    \I__397\ : Span12Mux_v
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__396\ : Odrv12
    port map (
            O => \N__4423\,
            I => \PIO_S0_c\
        );

    \I__395\ : ClkMux
    port map (
            O => \N__4420\,
            I => \N__4384\
        );

    \I__394\ : ClkMux
    port map (
            O => \N__4419\,
            I => \N__4384\
        );

    \I__393\ : ClkMux
    port map (
            O => \N__4418\,
            I => \N__4384\
        );

    \I__392\ : ClkMux
    port map (
            O => \N__4417\,
            I => \N__4384\
        );

    \I__391\ : ClkMux
    port map (
            O => \N__4416\,
            I => \N__4384\
        );

    \I__390\ : ClkMux
    port map (
            O => \N__4415\,
            I => \N__4384\
        );

    \I__389\ : ClkMux
    port map (
            O => \N__4414\,
            I => \N__4384\
        );

    \I__388\ : ClkMux
    port map (
            O => \N__4413\,
            I => \N__4384\
        );

    \I__387\ : ClkMux
    port map (
            O => \N__4412\,
            I => \N__4384\
        );

    \I__386\ : ClkMux
    port map (
            O => \N__4411\,
            I => \N__4384\
        );

    \I__385\ : ClkMux
    port map (
            O => \N__4410\,
            I => \N__4384\
        );

    \I__384\ : ClkMux
    port map (
            O => \N__4409\,
            I => \N__4384\
        );

    \I__383\ : GlobalMux
    port map (
            O => \N__4384\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            I => \N__4409\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__4415\
        );

    \INVU409_TRANSFER_ACK.TACK_OUTnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            I => \N__4413\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4411\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            I => \N__4410\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__4418\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__4417\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__4416\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            I => \N__4414\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            I => \N__4412\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            I => \N__4420\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            I => \N__4419\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_7C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            I => \N__10351\
        );

    \INVU409_AUTOCONFIG.ATA_BASE_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.ATA_BASE_2C_net\,
            I => \N__10357\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            I => \N__10348\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            I => \N__10359\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            I => \N__10349\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            I => \N__10352\
        );

    \INVU409_AUTOCONFIG.STATE_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_0C_net\,
            I => \N__10358\
        );

    \INVU409_AUTOCONFIG.LIDE_CONFC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            I => \N__10363\
        );

    \IN_MUX_bfv_14_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_5_0_\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_14_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_14_8_0_\
        );

    \IN_MUX_bfv_12_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10636\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_4_1_0_a2_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5564\,
            in2 => \_gnd_net_\,
            in3 => \N__6270\,
            lcout => \U409_AUTOCONFIG.N_214_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE10_2_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4532\,
            in1 => \N__4571\,
            in2 => \N__5802\,
            in3 => \N__5450\,
            lcout => \U409_AUTOCONFIG.ATA_BASE10Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_2_0__m2_0_123_i_i_a3_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5541\,
            in1 => \N__6244\,
            in2 => \N__5451\,
            in3 => \N__5693\,
            lcout => \U409_AUTOCONFIG.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__5694\,
            in2 => \_gnd_net_\,
            in3 => \N__5540\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_0_62_i_i_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_8_sqmuxa_i_o2_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000111111"
        )
    port map (
            in0 => \N__4479\,
            in1 => \N__5814\,
            in2 => \N__5712\,
            in3 => \N__5433\,
            lcout => \U409_AUTOCONFIG.N_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_2_0_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4588\,
            in1 => \N__5432\,
            in2 => \_gnd_net_\,
            in3 => \N__4533\,
            lcout => \U409_AUTOCONFIG.N_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_2_0_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4544\,
            in1 => \N__5788\,
            in2 => \N__4583\,
            in3 => \N__5466\,
            lcout => \U409_AUTOCONFIG.N_67\,
            ltout => \U409_AUTOCONFIG.N_67_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_1_LC_3_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__6294\,
            in1 => \N__10809\,
            in2 => \N__4483\,
            in3 => \N__5578\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_0_LC_3_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4543\,
            in2 => \_gnd_net_\,
            in3 => \N__4572\,
            lcout => \U409_AUTOCONFIG.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_2_LC_3_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__4545\,
            in2 => \N__4480\,
            in3 => \N__4576\,
            lcout => \U409_AUTOCONFIG.N_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_18_0_LC_3_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5579\,
            in1 => \N__6295\,
            in2 => \N__4584\,
            in3 => \N__5467\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.un1_A_18Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_18_LC_3_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5727\,
            in1 => \N__4546\,
            in2 => \N__4507\,
            in3 => \N__5789\,
            lcout => \U409_AUTOCONFIG.un1_AZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_4_0_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010101"
        )
    port map (
            in0 => \N__5816\,
            in1 => \N__6246\,
            in2 => \N__5464\,
            in3 => \N__5696\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_0_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__10832\,
            in1 => \N__4659\,
            in2 => \N__4504\,
            in3 => \N__5542\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_3_0_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5543\,
            in1 => \N__6245\,
            in2 => \_gnd_net_\,
            in3 => \N__5695\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a3_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010001000"
        )
    port map (
            in0 => \N__5115\,
            in1 => \N__4501\,
            in2 => \N__4495\,
            in3 => \N__5815\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_18_3_0_a2_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5697\,
            lcout => \U409_AUTOCONFIG.N_196_1\,
            ltout => \U409_AUTOCONFIG.N_196_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__6247\,
            in1 => \N__5455\,
            in2 => \N__4492\,
            in3 => \N__4489\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_3_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6074\,
            in1 => \N__10833\,
            in2 => \_gnd_net_\,
            in3 => \N__6026\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_5_LC_3_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6507\,
            in1 => \N__5279\,
            in2 => \N__5242\,
            in3 => \N__5341\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_3_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6607\,
            in1 => \N__4627\,
            in2 => \N__4621\,
            in3 => \N__5978\,
            lcout => \U409_ADDRESS_DECODE_Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8017\,
            in1 => \N__7489\,
            in2 => \_gnd_net_\,
            in3 => \N__7822\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__4998\,
            in1 => \N__4974\,
            in2 => \N__6406\,
            in3 => \N__6160\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9736\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4975\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9736\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5922\,
            in2 => \_gnd_net_\,
            in3 => \N__6782\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__9736\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0EA21_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5577\,
            in1 => \N__6154\,
            in2 => \N__5734\,
            in3 => \N__4618\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.ATA_BASE10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIH7AQ2_0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000000000"
        )
    port map (
            in0 => \N__4997\,
            in1 => \N__6372\,
            in2 => \N__4606\,
            in3 => \N__4966\,
            lcout => \U409_AUTOCONFIG.un1_STATE_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNISS061_3_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111100000"
        )
    port map (
            in0 => \N__5923\,
            in1 => \N__4732\,
            in2 => \N__6170\,
            in3 => \N__5089\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_a4_0_2_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7862\,
            in1 => \N__8215\,
            in2 => \_gnd_net_\,
            in3 => \N__8004\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.g0_i_a4_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_0_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__8522\,
            in1 => \N__7450\,
            in2 => \N__4738\,
            in3 => \N__5188\,
            lcout => \U409_ADDRESS_DECODE.g0_i_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10822\,
            in1 => \N__4973\,
            in2 => \N__4717\,
            in3 => \N__5182\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_3_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000100000"
        )
    port map (
            in0 => \N__4644\,
            in1 => \N__5580\,
            in2 => \N__6297\,
            in3 => \N__5728\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__10825\,
            in1 => \N__4728\,
            in2 => \N__4735\,
            in3 => \N__4798\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNIJJLA1_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6396\,
            in1 => \N__4965\,
            in2 => \N__4713\,
            in3 => \N__5181\,
            lcout => \U409_AUTOCONFIG.N_59_1\,
            ltout => \U409_AUTOCONFIG.N_59_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI777K2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__10823\,
            in1 => \N__4678\,
            in2 => \N__4666\,
            in3 => \N__4663\,
            lcout => \U409_AUTOCONFIG.AC_START_RNI777KZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__4770\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4633\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101010001000"
        )
    port map (
            in0 => \N__10824\,
            in1 => \N__5898\,
            in2 => \N__4648\,
            in3 => \N__4797\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_1_2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__4645\,
            in1 => \N__5581\,
            in2 => \N__6298\,
            in3 => \N__5729\,
            lcout => \U409_AUTOCONFIG.N_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000101"
        )
    port map (
            in0 => \N__4819\,
            in1 => \N__5031\,
            in2 => \N__4810\,
            in3 => \N__4783\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_6_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__7661\,
            in2 => \N__7780\,
            in3 => \N__7556\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI9THQ1_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10836\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4796\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa\,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_8_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__4777\,
            in1 => \N__4756\,
            in2 => \N__4744\,
            in3 => \N__5061\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5560\,
            in1 => \N__5701\,
            in2 => \N__6296\,
            in3 => \N__5448\,
            lcout => \U409_AUTOCONFIG.N_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_4_0_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7973\,
            in1 => \N__7414\,
            in2 => \N__8237\,
            in3 => \N__8488\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_1_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010001"
        )
    port map (
            in0 => \N__5733\,
            in1 => \N__5818\,
            in2 => \_gnd_net_\,
            in3 => \N__5465\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_7_94_i_i_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000110000"
        )
    port map (
            in0 => \N__5610\,
            in1 => \N__5559\,
            in2 => \N__4741\,
            in3 => \N__6233\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTc_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6619\,
            in1 => \N__6528\,
            in2 => \N__5293\,
            in3 => \N__5338\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5239\,
            in2 => \N__4939\,
            in3 => \N__6081\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4936\,
            in1 => \N__6032\,
            in2 => \_gnd_net_\,
            in3 => \N__5991\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4927\,
            in1 => \_gnd_net_\,
            in2 => \N__4921\,
            in3 => \N__4879\,
            lcout => \AUTOVECTOR\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6564\,
            in1 => \N__4918\,
            in2 => \N__4900\,
            in3 => \N__10840\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8418\,
            in1 => \N__8536\,
            in2 => \N__8236\,
            in3 => \N__7540\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4873\,
            in1 => \N__7770\,
            in2 => \N__4867\,
            in3 => \N__7621\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => \AUTOCONFIG_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4864\,
            in3 => \N__6401\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9919\,
            lcout => \un1_AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7267\,
            in1 => \N__6778\,
            in2 => \N__6892\,
            in3 => \N__5844\,
            lcout => \BRIDGE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.ATA_BASE_5_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7265\,
            in1 => \N__6803\,
            in2 => \N__6891\,
            in3 => \N__6659\,
            lcout => \ATA_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6777\,
            in2 => \_gnd_net_\,
            in3 => \N__6710\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.ATA_BASE_4_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7264\,
            in1 => \N__6802\,
            in2 => \N__6930\,
            in3 => \N__8096\,
            lcout => \ATA_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__6108\,
            in1 => \N__7266\,
            in2 => \N__6786\,
            in3 => \N__6926\,
            lcout => \BRIDGE_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__6850\,
            in2 => \N__7277\,
            in3 => \N__5829\,
            lcout => \BRIDGE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_1C_net\,
            ce => 'H',
            sr => \N__9735\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__5035\,
            in1 => \N__5924\,
            in2 => \N__5158\,
            in3 => \N__6159\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_a4_1_3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7451\,
            in1 => \N__8542\,
            in2 => \N__7877\,
            in3 => \N__8222\,
            lcout => \U409_ADDRESS_DECODE.g0_i_a4_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_12_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8388\,
            in1 => \N__7869\,
            in2 => \N__7486\,
            in3 => \N__8033\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.G_14_0_a7_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_10_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8543\,
            in2 => \N__5002\,
            in3 => \N__8223\,
            lcout => \U409_TRANSFER_ACK.N_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI25A42_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4999\,
            in1 => \N__4967\,
            in2 => \N__6387\,
            in3 => \N__6158\,
            lcout => \U409_AUTOCONFIG.BRIDGE_BASE_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_a4_1_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5194\,
            in1 => \N__8389\,
            in2 => \_gnd_net_\,
            in3 => \N__8010\,
            lcout => \U409_ADDRESS_DECODE.g0_i_a4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_1_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__7040\,
            in1 => \N__9291\,
            in2 => \_gnd_net_\,
            in3 => \N__7109\,
            lcout => \U409_ADDRESS_DECODE_ROMEN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__9929\,
            in1 => \N__9475\,
            in2 => \N__10808\,
            in3 => \N__6717\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10350\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__5170\,
            in1 => \N__5151\,
            in2 => \N__5362\,
            in3 => \N__5101\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9728\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101011100000010"
        )
    port map (
            in0 => \N__5102\,
            in1 => \N__5140\,
            in2 => \N__5134\,
            in3 => \N__5070\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9728\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010111001100"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__5883\,
            in2 => \N__5746\,
            in3 => \N__5103\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9728\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__5104\,
            in1 => \N__5641\,
            in2 => \N__5088\,
            in3 => \N__5745\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => 'H',
            sr => \N__9728\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100100"
        )
    port map (
            in0 => \N__6177\,
            in1 => \N__5071\,
            in2 => \N__5935\,
            in3 => \N__5062\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIQQ061_2_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__5934\,
            in1 => \N__5899\,
            in2 => \N__5887\,
            in3 => \N__6178\,
            lcout => \U409_AUTOCONFIG_D_OUT_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_0_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__5278\,
            in1 => \N__5334\,
            in2 => \N__5851\,
            in3 => \N__5833\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_0_3_144_i_i_a2_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5555\,
            in1 => \N__5810\,
            in2 => \N__6299\,
            in3 => \N__5702\,
            lcout => \U409_AUTOCONFIG.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_3_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6288\,
            in1 => \N__5449\,
            in2 => \N__5576\,
            in3 => \N__5703\,
            lcout => \U409_AUTOCONFIG.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5635\,
            in1 => \N__5611\,
            in2 => \N__5575\,
            in3 => \N__5431\,
            lcout => \U409_AUTOCONFIG.N_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6088\,
            in1 => \N__6621\,
            in2 => \N__5992\,
            in3 => \N__6036\,
            lcout => \U409_ADDRESS_DECODE.g2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_0_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5339\,
            in1 => \N__5291\,
            in2 => \N__10834\,
            in3 => \N__5240\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.g2_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_9_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__5944\,
            in2 => \N__5344\,
            in3 => \N__6716\,
            lcout => \U409_ADDRESS_DECODE.g2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_6_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5340\,
            in1 => \N__5292\,
            in2 => \N__10835\,
            in3 => \N__5241\,
            lcout => \U409_ADDRESS_DECODE_g2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_5_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6620\,
            in1 => \N__6087\,
            in2 => \N__6037\,
            in3 => \N__5987\,
            lcout => \U409_ADDRESS_DECODE.g2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_4_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7013\,
            in1 => \N__7086\,
            in2 => \_gnd_net_\,
            in3 => \N__6529\,
            lcout => \U409_ADDRESS_DECODE.g2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_1_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__8537\,
            in1 => \N__6658\,
            in2 => \N__8252\,
            in3 => \N__8092\,
            lcout => \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_9_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7824\,
            in1 => \N__7491\,
            in2 => \N__8253\,
            in3 => \N__8538\,
            lcout => \U409_TRANSFER_ACK.G_14_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_10_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__7823\,
            in1 => \N__7185\,
            in2 => \N__7779\,
            in3 => \N__6946\,
            lcout => \U409_ADDRESS_DECODE.g2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_o4_1_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__7343\,
            in1 => \N__7658\,
            in2 => \N__7596\,
            in3 => \N__7552\,
            lcout => \U409_ADDRESS_DECODE.g0_i_o4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_6_0_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__7659\,
            in1 => \N__7588\,
            in2 => \N__7558\,
            in3 => \N__7342\,
            lcout => \U409_ADDRESS_DECODE.un1_Z2_SPACE_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000100"
        )
    port map (
            in0 => \N__8119\,
            in1 => \N__8419\,
            in2 => \N__8028\,
            in3 => \N__6698\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7481\,
            in2 => \N__5938\,
            in3 => \N__7318\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_Z2_SPACE_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6421\,
            in1 => \N__6415\,
            in2 => \N__6409\,
            in3 => \N__7570\,
            lcout => \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.un1_Z2_SPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_ROM_EN_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__6400\,
            in1 => \N__9492\,
            in2 => \N__6328\,
            in3 => \N__10014\,
            lcout => \U409_ADDRESS_DECODE_ATA_ROM_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10356\,
            ce => 'H',
            sr => \N__9733\
        );

    \U409_ADDRESS_DECODE.g2_11_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__7490\,
            in1 => \N__7323\,
            in2 => \N__8040\,
            in3 => \N__8126\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.g2Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITNPB5_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010101010101"
        )
    port map (
            in0 => \N__10015\,
            in1 => \N__6325\,
            in2 => \N__6316\,
            in3 => \N__6313\,
            lcout => \U409_ADDRESS_DECODE_ATA_ROM_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI0FVT2_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__6120\,
            in1 => \N__6301\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.STATE_RNI0FVT2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9A3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6300\,
            in1 => \N__6176\,
            in2 => \_gnd_net_\,
            in3 => \N__6121\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIHQ9AZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8626\,
            in2 => \_gnd_net_\,
            in3 => \N__8753\,
            lcout => \U409_TRANSFER_ACK.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_2_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000010001"
        )
    port map (
            in0 => \N__6715\,
            in1 => \N__6527\,
            in2 => \_gnd_net_\,
            in3 => \N__6109\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_4_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__7041\,
            in1 => \N__7110\,
            in2 => \N__6091\,
            in3 => \N__10776\,
            lcout => \U409_ADDRESS_DECODE.un1_BRIDGE_ENnZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_8_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__8532\,
            in1 => \N__6451\,
            in2 => \N__6670\,
            in3 => \N__6714\,
            lcout => \U409_TRANSFER_ACK.G_14_0_o7_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g0_i_o4_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__6669\,
            in1 => \N__8098\,
            in2 => \N__8241\,
            in3 => \N__8531\,
            lcout => \U409_ADDRESS_DECODE.g0_i_o4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BRIDGE_ENn_i_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110111111"
        )
    port map (
            in0 => \N__6748\,
            in1 => \N__6640\,
            in2 => \N__6634\,
            in3 => \N__6625\,
            lcout => \U409_ADDRESS_DECODE_un1_BRIDGE_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6565\,
            in1 => \N__8505\,
            in2 => \_gnd_net_\,
            in3 => \N__8221\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6541\,
            in1 => \N__7487\,
            in2 => \N__6544\,
            in3 => \N__9276\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7030\,
            in1 => \N__7099\,
            in2 => \_gnd_net_\,
            in3 => \N__8018\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.g2_7_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001000"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__6535\,
            in2 => \N__7085\,
            in3 => \N__6517\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE_g2_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_11_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__6460\,
            in1 => \_gnd_net_\,
            in2 => \N__6454\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.G_14_0_o7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__9304\,
            in1 => \N__6967\,
            in2 => \N__7665\,
            in3 => \N__6955\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_3_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8251\,
            in1 => \N__8548\,
            in2 => \N__7870\,
            in3 => \N__7734\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6966\,
            in1 => \N__9303\,
            in2 => \N__6949\,
            in3 => \N__7654\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_Z2_SPACE_7_2_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__7735\,
            in1 => \N__7838\,
            in2 => \N__7186\,
            in3 => \N__6944\,
            lcout => \U409_ADDRESS_DECODE_un1_Z2_SPACE_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.ATA_BASE_2_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__6945\,
            in1 => \N__7278\,
            in2 => \N__6846\,
            in3 => \N__7240\,
            lcout => \ATA_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_2C_net\,
            ce => 'H',
            sr => \N__9734\
        );

    \U409_AUTOCONFIG.ATA_BASE_7_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__7217\,
            in1 => \N__6805\,
            in2 => \N__8127\,
            in3 => \N__7296\,
            lcout => \ATA_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_AUTOCONFIG.ATA_BASE_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7292\,
            in1 => \N__7234\,
            in2 => \N__6931\,
            in3 => \N__7344\,
            lcout => \ATA_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_AUTOCONFIG.ATA_BASE_1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__7293\,
            in1 => \N__7235\,
            in2 => \N__7597\,
            in3 => \N__6873\,
            lcout => \ATA_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_AUTOCONFIG.ATA_BASE_6_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__6836\,
            in1 => \N__6804\,
            in2 => \N__7324\,
            in3 => \N__7295\,
            lcout => \ATA_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__7218\,
            in1 => \N__7297\,
            in2 => \N__6747\,
            in3 => \N__6787\,
            lcout => \BRIDGE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_AUTOCONFIG.ATA_BASE_3_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7294\,
            in1 => \N__7236\,
            in2 => \N__7219\,
            in3 => \N__7184\,
            lcout => \ATA_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.ATA_BASE_7C_net\,
            ce => 'H',
            sr => \N__9730\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8627\,
            in2 => \_gnd_net_\,
            in3 => \N__8754\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__9729\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__7132\,
            in1 => \N__8062\,
            in2 => \N__7165\,
            in3 => \N__8056\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__9729\
        );

    \U409_ADDRESS_DECODE.ATA_ROM_EN_RNITAAO4_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010101"
        )
    port map (
            in0 => \N__7156\,
            in1 => \N__7147\,
            in2 => \N__10034\,
            in3 => \N__7138\,
            lcout => \U409_ADDRESS_DECODE_ATA_ROM_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000010100"
        )
    port map (
            in0 => \N__8590\,
            in1 => \N__7125\,
            in2 => \N__8668\,
            in3 => \N__8572\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__9726\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__8663\,
            in1 => \N__8554\,
            in2 => \N__7126\,
            in3 => \N__8795\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__9726\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_2_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__7111\,
            in1 => \N__7488\,
            in2 => \N__7042\,
            in3 => \N__7969\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011111111"
        )
    port map (
            in0 => \N__8217\,
            in1 => \N__7879\,
            in2 => \N__7778\,
            in3 => \N__7687\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un2_REGSPACEn_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un2_REGSPACEn_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__8545\,
            in1 => \N__7693\,
            in2 => \N__7882\,
            in3 => \N__7699\,
            lcout => \U409_ADDRESS_DECODE_un2_REGSPACEn_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.REG_SPACE_2_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8216\,
            in1 => \N__7878\,
            in2 => \N__7777\,
            in3 => \N__7666\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_4_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8029\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7461\,
            lcout => \U409_ADDRESS_DECODE.REG_SPACE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.RAN_SPACE_0_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__7462\,
            in1 => \N__8030\,
            in2 => \_gnd_net_\,
            in3 => \N__8544\,
            lcout => \U409_ADDRESS_DECODE.RAN_SPACEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8041\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7492\,
            lcout => \U409_ADDRESS_DECODE.LOWROMZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_RNO_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__8925\,
            in1 => \N__8940\,
            in2 => \_gnd_net_\,
            in3 => \N__9498\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERc_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__8547\,
            in1 => \N__8434\,
            in2 => \N__8387\,
            in3 => \N__8304\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_4_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011111111"
        )
    port map (
            in0 => \N__7660\,
            in1 => \N__7595\,
            in2 => \_gnd_net_\,
            in3 => \N__7569\,
            lcout => \U409_TRANSFER_ACK.g0_0_0_o6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_6_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__7557\,
            in1 => \N__7482\,
            in2 => \N__7348\,
            in3 => \N__7322\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.G_14_0_o7_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_3_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__8068\,
            in1 => \_gnd_net_\,
            in2 => \N__8269\,
            in3 => \N__8266\,
            lcout => \U409_TRANSFER_ACK.G_14_0_o7_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_7_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__8032\,
            in1 => \N__8254\,
            in2 => \N__8128\,
            in3 => \N__8097\,
            lcout => \U409_TRANSFER_ACK.G_14_0_o7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100010001"
        )
    port map (
            in0 => \N__8055\,
            in1 => \N__8589\,
            in2 => \N__8680\,
            in3 => \N__8571\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101011"
        )
    port map (
            in0 => \N__8750\,
            in1 => \N__8623\,
            in2 => \N__8667\,
            in3 => \N__8787\,
            lcout => \U409_TRANSFER_ACK.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_1_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8786\,
            in1 => \N__8657\,
            in2 => \N__8629\,
            in3 => \N__8749\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__8588\,
            in1 => \_gnd_net_\,
            in2 => \N__8044\,
            in3 => \N__8676\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__8625\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8662\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_5_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__8031\,
            in1 => \N__7909\,
            in2 => \N__7900\,
            in3 => \N__8788\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.G_14_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_2_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8624\,
            in1 => \N__8661\,
            in2 => \N__7885\,
            in3 => \N__8751\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.G_14_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__8698\,
            in1 => \N__10035\,
            in2 => \N__8689\,
            in3 => \N__8686\,
            lcout => \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_s_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__8420\,
            in1 => \N__9488\,
            in2 => \_gnd_net_\,
            in3 => \N__10388\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIAR8J_0_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8656\,
            in1 => \N__8752\,
            in2 => \N__8628\,
            in3 => \N__8789\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_3_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8575\,
            in3 => \N__8570\,
            lcout => \U409_TRANSFER_ACK.ROMENn_1_sqmuxa_0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__8546\,
            in1 => \N__8433\,
            in2 => \N__8377\,
            in3 => \N__8311\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9295\,
            in2 => \_gnd_net_\,
            in3 => \N__9315\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => \U409_ADDRESS_DECODE_un1_REGSPACEn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9947\,
            in1 => \N__8956\,
            in2 => \N__8293\,
            in3 => \N__9896\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__8902\,
            in1 => \N__8965\,
            in2 => \N__8881\,
            in3 => \N__10391\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9731\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__8971\,
            in1 => \N__10390\,
            in2 => \_gnd_net_\,
            in3 => \N__8964\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9731\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__10741\,
            in1 => \N__8952\,
            in2 => \N__8929\,
            in3 => \N__9499\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10752\,
            in1 => \N__9652\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNI7KT7_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8860\,
            in3 => \N__8709\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIBQIN_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8896\,
            in1 => \N__8877\,
            in2 => \N__8866\,
            in3 => \N__9510\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001010"
        )
    port map (
            in0 => \N__10751\,
            in1 => \N__9653\,
            in2 => \N__8863\,
            in3 => \N__9675\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111100001000"
        )
    port map (
            in0 => \N__10207\,
            in1 => \N__9688\,
            in2 => \N__10237\,
            in3 => \N__8859\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__8817\,
            in1 => \N__8845\,
            in2 => \N__8806\,
            in3 => \N__8839\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100100000"
        )
    port map (
            in0 => \N__8802\,
            in1 => \N__8761\,
            in2 => \N__8719\,
            in3 => \N__8710\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10431\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000001110001"
        )
    port map (
            in0 => \N__9655\,
            in1 => \N__9676\,
            in2 => \N__9848\,
            in3 => \N__9628\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9550\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__9727\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI1CKM1_7_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9022\,
            in1 => \N__9046\,
            in2 => \N__9127\,
            in3 => \N__8987\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_4_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__9412\,
            in1 => \N__10105\,
            in2 => \N__8992\,
            in3 => \N__9106\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__10106\,
            in1 => \N__9025\,
            in2 => \N__10156\,
            in3 => \N__10134\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10080\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__9126\,
            in1 => \N__9004\,
            in2 => \N__10138\,
            in3 => \N__8989\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10080\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIO2KM1_3_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__9023\,
            in1 => \N__9413\,
            in2 => \N__9052\,
            in3 => \N__10104\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_7_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__9125\,
            in1 => \N__8988\,
            in2 => \N__8974\,
            in3 => \N__9105\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_7_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__9493\,
            in1 => \N__10387\,
            in2 => \N__9133\,
            in3 => \N__9527\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9124\,
            in2 => \N__9130\,
            in3 => \N__9003\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10080\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__9416\,
            in1 => \N__9094\,
            in2 => \_gnd_net_\,
            in3 => \N__10132\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10076\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__9093\,
            in1 => \_gnd_net_\,
            in2 => \N__9076\,
            in3 => \N__9418\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10076\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9090\,
            in2 => \_gnd_net_\,
            in3 => \N__9064\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__9092\,
            in1 => \_gnd_net_\,
            in2 => \N__9075\,
            in3 => \N__9415\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__9051\,
            in1 => \_gnd_net_\,
            in2 => \N__9097\,
            in3 => \N__10131\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10076\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9091\,
            in1 => \N__9414\,
            in2 => \N__9074\,
            in3 => \N__9050\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10111\,
            in2 => \N__9028\,
            in3 => \N__9024\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__9497\,
            in1 => \N__9417\,
            in2 => \N__10393\,
            in3 => \N__9529\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10076\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__9391\,
            in1 => \N__9354\,
            in2 => \N__9385\,
            in3 => \N__10767\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_DATA_BUFFERS.un1_BUFENn_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__9325\,
            in1 => \N__9297\,
            in2 => \N__9361\,
            in3 => \N__9948\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9296\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10695\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9970\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9220\,
            in3 => \N__9217\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9172\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10270\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10724\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9969\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_1C_net\,
            ce => 'H',
            sr => \N__9732\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__10283\,
            in1 => \N__10268\,
            in2 => \N__10202\,
            in3 => \N__9687\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__10739\,
            in1 => \N__10230\,
            in2 => \N__9697\,
            in3 => \N__9694\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111100010000"
        )
    port map (
            in0 => \N__10284\,
            in1 => \N__10267\,
            in2 => \N__10203\,
            in3 => \N__10248\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9549\,
            in1 => \N__10389\,
            in2 => \_gnd_net_\,
            in3 => \N__9562\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100111"
        )
    port map (
            in0 => \N__9673\,
            in1 => \N__9575\,
            in2 => \N__9654\,
            in3 => \N__9627\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000101110"
        )
    port map (
            in0 => \N__9576\,
            in1 => \N__10740\,
            in2 => \N__9616\,
            in3 => \_gnd_net_\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_OUTnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9561\,
            in2 => \_gnd_net_\,
            in3 => \N__9548\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__9511\,
            in1 => \N__9535\,
            in2 => \_gnd_net_\,
            in3 => \N__9528\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10081\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__10155\,
            in1 => \N__10110\,
            in2 => \_gnd_net_\,
            in3 => \N__10133\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10081\
        );

    \U409_ADDRESS_DECODE.ATA_ROM_EN_RNIBHHS6_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10048\,
            in2 => \_gnd_net_\,
            in3 => \N__10036\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10884\,
            in2 => \_gnd_net_\,
            in3 => \N__10537\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10480\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10556\,
            in2 => \_gnd_net_\,
            in3 => \N__10577\,
            lcout => \U409_CIA.CLK_CIA6_4\,
            ltout => \U409_CIA.CLK_CIA6_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__10591\,
            in1 => \N__10462\,
            in2 => \N__9976\,
            in3 => \N__10535\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__10536\,
            in1 => \N__9901\,
            in2 => \N__9973\,
            in3 => \N__9962\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10883\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10478\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNI1IRLB_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__9949\,
            in1 => \N__9897\,
            in2 => \_gnd_net_\,
            in3 => \N__9855\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10392\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__10285\,
            in1 => \N__10269\,
            in2 => \N__10201\,
            in3 => \N__10249\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__10714\,
            in1 => \N__10229\,
            in2 => \N__10210\,
            in3 => \N__10191\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10532\,
            in2 => \N__10885\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10924\,
            in2 => \_gnd_net_\,
            in3 => \N__10168\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__10479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10942\,
            in2 => \_gnd_net_\,
            in3 => \N__10165\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10459\,
            in2 => \_gnd_net_\,
            in3 => \N__10162\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__10479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10903\,
            in2 => \_gnd_net_\,
            in3 => \N__10159\,
            lcout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10579\,
            in2 => \_gnd_net_\,
            in3 => \N__10597\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__10479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10560\,
            in2 => \_gnd_net_\,
            in3 => \N__10594\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10479\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__10943\,
            in1 => \N__10925\,
            in2 => \N__10908\,
            in3 => \N__10880\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10852\,
            in1 => \N__10507\,
            in2 => \N__10501\,
            in3 => \N__10585\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10578\,
            in1 => \N__10882\,
            in2 => \N__10561\,
            in3 => \N__10534\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001101100"
        )
    port map (
            in0 => \N__10399\,
            in1 => \N__10417\,
            in2 => \N__10540\,
            in3 => \N__10907\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNI9DRM_4_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10460\,
            in2 => \_gnd_net_\,
            in3 => \N__10533\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__10497\,
            in1 => \N__10851\,
            in2 => \N__10489\,
            in3 => \N__10486\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10477\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011000"
        )
    port map (
            in0 => \N__10945\,
            in1 => \N__10461\,
            in2 => \N__10424\,
            in3 => \N__10927\,
            lcout => \U409_CIA.CLK_CIA_r_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10944\,
            in1 => \N__10926\,
            in2 => \N__10909\,
            in3 => \N__10881\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11193\,
            in2 => \_gnd_net_\,
            in3 => \N__11214\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__11043\,
            in1 => \N__10997\,
            in2 => \N__11461\,
            in3 => \N__11069\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__11042\,
            in1 => \N__11125\,
            in2 => \N__11002\,
            in3 => \N__11068\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNINQJI1_4_LC_13_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__11098\,
            in1 => \N__11137\,
            in2 => \N__11116\,
            in3 => \N__11473\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__11497\,
            in1 => \N__11045\,
            in2 => \N__10624\,
            in3 => \N__10998\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__10996\,
            in1 => \N__10608\,
            in2 => \N__11077\,
            in3 => \N__11044\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11075\,
            in1 => \N__10995\,
            in2 => \N__11047\,
            in3 => \N__11662\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIA84S_11_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11410\,
            in1 => \N__11152\,
            in2 => \N__11170\,
            in3 => \N__11395\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11074\,
            in1 => \N__10994\,
            in2 => \N__11046\,
            in3 => \N__11350\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIRP4S_14_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__11674\,
            in1 => \N__11449\,
            in2 => \N__11365\,
            in3 => \N__11488\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__11073\,
            in1 => \N__10993\,
            in2 => \N__11080\,
            in3 => \N__11192\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__10992\,
            in1 => \N__11076\,
            in2 => \N__11437\,
            in3 => \N__11041\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11847\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDAFF_10_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11380\,
            in1 => \N__11425\,
            in2 => \_gnd_net_\,
            in3 => \N__11191\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIVPLP1_16_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__11215\,
            in1 => \N__11649\,
            in2 => \N__11011\,
            in3 => \N__11008\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__11290\,
            in1 => \N__11323\,
            in2 => \N__11536\,
            in3 => \N__11248\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__11247\,
            in1 => \N__10956\,
            in2 => \N__11329\,
            in3 => \N__11292\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__11291\,
            in1 => \N__11324\,
            in2 => \N__11509\,
            in3 => \N__11249\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNI3J3V_10_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11770\,
            in1 => \N__11596\,
            in2 => \N__11638\,
            in3 => \N__11731\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11322\,
            in1 => \N__11289\,
            in2 => \N__11258\,
            in3 => \N__11740\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11637\,
            in2 => \_gnd_net_\,
            in3 => \N__11619\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11849\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11286\,
            in1 => \N__11320\,
            in2 => \N__11260\,
            in3 => \N__11704\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIJAR11_3_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11524\,
            in1 => \N__11581\,
            in2 => \N__11551\,
            in3 => \N__11791\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11287\,
            in1 => \N__11257\,
            in2 => \N__11086\,
            in3 => \N__11878\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIDMCS_11_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11695\,
            in1 => \N__11716\,
            in2 => \N__11755\,
            in3 => \N__11890\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11288\,
            in1 => \N__11321\,
            in2 => \N__11083\,
            in3 => \N__11779\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIG9CP_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11821\,
            in1 => \N__11566\,
            in2 => \_gnd_net_\,
            in3 => \N__11617\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNI02282_16_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__11865\,
            in1 => \N__11341\,
            in2 => \N__11335\,
            in3 => \N__11806\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__11319\,
            in1 => \N__11253\,
            in2 => \N__11332\,
            in3 => \N__11618\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11851\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__11328\,
            in1 => \N__11293\,
            in2 => \N__11259\,
            in3 => \N__11683\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11853\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11210\,
            in2 => \N__11194\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_5_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11166\,
            in2 => \_gnd_net_\,
            in3 => \N__11155\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__11848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11151\,
            in2 => \_gnd_net_\,
            in3 => \N__11140\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__11848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_14_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11136\,
            in2 => \_gnd_net_\,
            in3 => \N__11119\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11112\,
            in2 => \_gnd_net_\,
            in3 => \N__11101\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__11848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_14_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11097\,
            in2 => \_gnd_net_\,
            in3 => \N__11491\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_14_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11487\,
            in2 => \_gnd_net_\,
            in3 => \N__11476\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__11848\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11472\,
            in2 => \_gnd_net_\,
            in3 => \N__11452\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11448\,
            in2 => \_gnd_net_\,
            in3 => \N__11428\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11424\,
            in2 => \_gnd_net_\,
            in3 => \N__11413\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__11850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11409\,
            in2 => \_gnd_net_\,
            in3 => \N__11398\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__11850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11394\,
            in2 => \_gnd_net_\,
            in3 => \N__11383\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__11850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11379\,
            in2 => \_gnd_net_\,
            in3 => \N__11368\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__11850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11361\,
            in2 => \_gnd_net_\,
            in3 => \N__11344\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11673\,
            in2 => \_gnd_net_\,
            in3 => \N__11656\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11650\,
            in2 => \_gnd_net_\,
            in3 => \N__11653\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11850\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11633\,
            in2 => \N__11620\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11595\,
            in2 => \_gnd_net_\,
            in3 => \N__11584\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__11852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11580\,
            in2 => \_gnd_net_\,
            in3 => \N__11569\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__11852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11565\,
            in2 => \_gnd_net_\,
            in3 => \N__11554\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__11852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11547\,
            in2 => \_gnd_net_\,
            in3 => \N__11527\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11520\,
            in2 => \_gnd_net_\,
            in3 => \N__11500\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11820\,
            in2 => \_gnd_net_\,
            in3 => \N__11809\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__11852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11805\,
            in2 => \_gnd_net_\,
            in3 => \N__11794\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__11852\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11790\,
            in2 => \_gnd_net_\,
            in3 => \N__11773\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_8_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11769\,
            in2 => \_gnd_net_\,
            in3 => \N__11758\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__11854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11751\,
            in2 => \_gnd_net_\,
            in3 => \N__11734\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11730\,
            in2 => \_gnd_net_\,
            in3 => \N__11719\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__11854\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11715\,
            in2 => \_gnd_net_\,
            in3 => \N__11698\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11694\,
            in2 => \_gnd_net_\,
            in3 => \N__11677\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11889\,
            in2 => \_gnd_net_\,
            in3 => \N__11872\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11866\,
            in2 => \_gnd_net_\,
            in3 => \N__11869\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11854\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 25 2025 21:58:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    TICK50 : out std_logic;
    nROMEN : out std_logic;
    nCIACS1 : out std_logic;
    TICK60 : out std_logic;
    CLKCIA : out std_logic;
    CLK6 : in std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    TSn : in std_logic;
    nBUFEN : out std_logic;
    nREGSPACE : out std_logic;
    nRAMSPACE : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    TACKn : inout std_logic;
    nCIACS0 : out std_logic;
    PORTSIZE : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__6546\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6354\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6291\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6125\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5798\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5790\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5769\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5580\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4652\ : std_logic;
signal \N__4649\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4464\ : std_logic;
signal \N__4461\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4428\ : std_logic;
signal \N__4425\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4389\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4269\ : std_logic;
signal \N__4266\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3927\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3918\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3843\ : std_logic;
signal \N__3840\ : std_logic;
signal \N__3837\ : std_logic;
signal \N__3834\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3747\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3723\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3483\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3450\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3254\ : std_logic;
signal \N__3251\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3200\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3176\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3091\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2890\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2877\ : std_logic;
signal \N__2872\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2866\ : std_logic;
signal \N__2863\ : std_logic;
signal \N__2860\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2841\ : std_logic;
signal \N__2838\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2792\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2763\ : std_logic;
signal \N__2760\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2714\ : std_logic;
signal \N__2711\ : std_logic;
signal \N__2708\ : std_logic;
signal \N__2707\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2699\ : std_logic;
signal \N__2696\ : std_logic;
signal \N__2693\ : std_logic;
signal \N__2690\ : std_logic;
signal \N__2687\ : std_logic;
signal \N__2684\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2676\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2663\ : std_logic;
signal \N__2660\ : std_logic;
signal \N__2657\ : std_logic;
signal \N__2654\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2649\ : std_logic;
signal \N__2646\ : std_logic;
signal \N__2639\ : std_logic;
signal \N__2636\ : std_logic;
signal \N__2633\ : std_logic;
signal \N__2630\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2597\ : std_logic;
signal \N__2594\ : std_logic;
signal \N__2591\ : std_logic;
signal \N__2588\ : std_logic;
signal \N__2585\ : std_logic;
signal \N__2582\ : std_logic;
signal \N__2579\ : std_logic;
signal \N__2576\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2570\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2555\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2551\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2540\ : std_logic;
signal \N__2537\ : std_logic;
signal \N__2534\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2528\ : std_logic;
signal \N__2525\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2519\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2504\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2502\ : std_logic;
signal \N__2501\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2499\ : std_logic;
signal \N__2498\ : std_logic;
signal \N__2497\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2474\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U409_CIA.g0Z0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_CIA.g0Z0Z_10\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\ : std_logic;
signal \U409_CIA.g0Z0Z_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_CIA.g0Z0Z_11\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_6\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACEm_3\ : std_logic;
signal \A_c_19\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nREGSPACE_i\ : std_logic;
signal \bfn_11_5_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_11_6_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.m9_am_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.i6_mux_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_105_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.m9_bm\ : std_logic;
signal \U409_TRANSFER_ACK.N_4\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_23\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_ADDRESS_DECODE.LOWROMZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.HIROMZ0\ : std_logic;
signal \ROMENm_i\ : std_logic;
signal \AUTOVECTORm\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \ROMENm\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS0_i\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nCIACS1_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \CIA_ENABLEm\ : std_logic;
signal \U409_CIA.N_9_cascade_\ : std_logic;
signal \U409_CIA.g0Z0Z_14\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_CIA.g0Z0Z_13\ : std_logic;
signal \U409_CIA.CIA_HOLDZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_105\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \bfn_13_7_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\ : std_logic;
signal \U409_CIA.N_20_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CLKCIAZ0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \CLKCIA_c\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CLKCIA6_0_a2_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CLKCIA8_0_a2_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACEZ0\ : std_logic;
signal \OVL_c\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_EN_iC_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \nBUFEN_c\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \TACK_EN_i\ : std_logic;
signal \N_365_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \CLKCIA_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \nCIACS0_wire\ : std_logic;
signal \nCIACS1_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \nRAMSPACE_wire\ : std_logic;
signal \nROMEN_wire\ : std_logic;
signal \nBUFEN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \nREGSPACE_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \TT_wire\ <= TT;
    CLKCIA <= \CLKCIA_wire\;
    \A_wire\ <= A;
    nCIACS0 <= \nCIACS0_wire\;
    nCIACS1 <= \nCIACS1_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    nRAMSPACE <= \nRAMSPACE_wire\;
    nROMEN <= \nROMEN_wire\;
    nBUFEN <= \nBUFEN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    nREGSPACE <= \nREGSPACE_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TICK60 <= \TICK60_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__4118\,
            RESETB => \N__4040\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6544\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6546\,
            DIN => \N__6545\,
            DOUT => \N__6544\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6546\,
            PADOUT => \N__6545\,
            PADIN => \N__6544\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__6534\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6536\,
            DIN => \N__6535\,
            DOUT => \N__6534\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6536\,
            PADOUT => \N__6535\,
            PADIN => \N__6534\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6525\,
            DIN => \N__6524\,
            DOUT => \N__6523\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6525\,
            PADOUT => \N__6524\,
            PADIN => \N__6523\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKCIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6516\,
            DIN => \N__6515\,
            DOUT => \N__6514\,
            PACKAGEPIN => \CLKCIA_wire\
        );

    \CLKCIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6516\,
            PADOUT => \N__6515\,
            PADIN => \N__6514\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5417\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6507\,
            DIN => \N__6506\,
            DOUT => \N__6505\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6507\,
            PADOUT => \N__6506\,
            PADIN => \N__6505\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6498\,
            DIN => \N__6497\,
            DOUT => \N__6496\,
            PACKAGEPIN => \nCIACS0_wire\
        );

    \nCIACS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6498\,
            PADOUT => \N__6497\,
            PADIN => \N__6496\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4010\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nCIACS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6489\,
            DIN => \N__6488\,
            DOUT => \N__6487\,
            PACKAGEPIN => \nCIACS1_wire\
        );

    \nCIACS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6489\,
            PADOUT => \N__6488\,
            PADIN => \N__6487\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4628\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6480\,
            DIN => \N__6479\,
            DOUT => \N__6478\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6480\,
            PADOUT => \N__6479\,
            PADIN => \N__6478\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6471\,
            DIN => \N__6470\,
            DOUT => \N__6469\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6471\,
            PADOUT => \N__6470\,
            PADIN => \N__6469\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6462\,
            DIN => \N__6461\,
            DOUT => \N__6460\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6462\,
            PADOUT => \N__6461\,
            PADIN => \N__6460\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6453\,
            DIN => \N__6452\,
            DOUT => \N__6451\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__6453\,
            PADOUT => \N__6452\,
            PADIN => \N__6451\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5885\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__5555\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6444\,
            DIN => \N__6443\,
            DOUT => \N__6442\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6444\,
            PADOUT => \N__6443\,
            PADIN => \N__6442\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6435\,
            DIN => \N__6434\,
            DOUT => \N__6433\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6435\,
            PADOUT => \N__6434\,
            PADIN => \N__6433\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6426\,
            DIN => \N__6425\,
            DOUT => \N__6424\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6426\,
            PADOUT => \N__6425\,
            PADIN => \N__6424\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6417\,
            DIN => \N__6416\,
            DOUT => \N__6415\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6417\,
            PADOUT => \N__6416\,
            PADIN => \N__6415\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nRAMSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6408\,
            DIN => \N__6407\,
            DOUT => \N__6406\,
            PACKAGEPIN => \nRAMSPACE_wire\
        );

    \nRAMSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6408\,
            PADOUT => \N__6407\,
            PADIN => \N__6406\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4613\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nROMEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6399\,
            DIN => \N__6398\,
            DOUT => \N__6397\,
            PACKAGEPIN => \nROMEN_wire\
        );

    \nROMEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6399\,
            PADOUT => \N__6398\,
            PADIN => \N__6397\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6390\,
            DIN => \N__6389\,
            DOUT => \N__6388\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6390\,
            PADOUT => \N__6389\,
            PADIN => \N__6388\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6381\,
            DIN => \N__6380\,
            DOUT => \N__6379\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6381\,
            PADOUT => \N__6380\,
            PADIN => \N__6379\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nBUFEN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6372\,
            DIN => \N__6371\,
            DOUT => \N__6370\,
            PACKAGEPIN => \nBUFEN_wire\
        );

    \nBUFEN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6372\,
            PADOUT => \N__6371\,
            PADIN => \N__6370\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6363\,
            DIN => \N__6362\,
            DOUT => \N__6361\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6363\,
            PADOUT => \N__6362\,
            PADIN => \N__6361\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6354\,
            DIN => \N__6353\,
            DOUT => \N__6352\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6354\,
            PADOUT => \N__6353\,
            PADIN => \N__6352\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6345\,
            DIN => \N__6344\,
            DOUT => \N__6343\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6345\,
            PADOUT => \N__6344\,
            PADIN => \N__6343\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6336\,
            DIN => \N__6335\,
            DOUT => \N__6334\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6336\,
            PADOUT => \N__6335\,
            PADIN => \N__6334\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6327\,
            DIN => \N__6326\,
            DOUT => \N__6325\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6327\,
            PADOUT => \N__6326\,
            PADIN => \N__6325\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6318\,
            DIN => \N__6317\,
            DOUT => \N__6316\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6318\,
            PADOUT => \N__6317\,
            PADIN => \N__6316\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6309\,
            DIN => \N__6308\,
            DOUT => \N__6307\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6309\,
            PADOUT => \N__6308\,
            PADIN => \N__6307\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \nREGSPACE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6300\,
            DIN => \N__6299\,
            DOUT => \N__6298\,
            PACKAGEPIN => \nREGSPACE_wire\
        );

    \nREGSPACE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6300\,
            PADOUT => \N__6299\,
            PADIN => \N__6298\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3611\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6291\,
            DIN => \N__6290\,
            DOUT => \N__6289\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6291\,
            PADOUT => \N__6290\,
            PADIN => \N__6289\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3572\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6282\,
            DIN => \N__6281\,
            DOUT => \N__6280\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6282\,
            PADOUT => \N__6281\,
            PADIN => \N__6280\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6273\,
            DIN => \N__6272\,
            DOUT => \N__6271\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6273\,
            PADOUT => \N__6272\,
            PADIN => \N__6271\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6264\,
            DIN => \N__6263\,
            DOUT => \N__6262\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6264\,
            PADOUT => \N__6263\,
            PADIN => \N__6262\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6255\,
            DIN => \N__6254\,
            DOUT => \N__6253\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6255\,
            PADOUT => \N__6254\,
            PADIN => \N__6253\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6246\,
            DIN => \N__6245\,
            DOUT => \N__6244\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6246\,
            PADOUT => \N__6245\,
            PADIN => \N__6244\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6237\,
            DIN => \N__6236\,
            DOUT => \N__6235\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6237\,
            PADOUT => \N__6236\,
            PADIN => \N__6235\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4595\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6228\,
            DIN => \N__6227\,
            DOUT => \N__6226\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6228\,
            PADOUT => \N__6227\,
            PADIN => \N__6226\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__6219\,
            DIN => \N__6218\,
            DOUT => \N__6217\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6219\,
            PADOUT => \N__6218\,
            PADIN => \N__6217\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__6200\,
            I => \N__6195\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6188\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6188\
        );

    \I__1454\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6188\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__6188\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6176\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6184\,
            I => \N__6176\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6183\,
            I => \N__6176\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6176\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6173\,
            I => \N__6169\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6172\,
            I => \N__6166\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6169\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__6166\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\
        );

    \I__1444\ : CEMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1442\ : Odrv4
    port map (
            O => \N__6155\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6148\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__6151\,
            I => \N__6144\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6148\,
            I => \N__6141\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6138\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6144\,
            I => \N__6135\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__6141\,
            I => \N__6132\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6138\,
            I => \N__6127\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6135\,
            I => \N__6127\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__6132\,
            I => \N__6120\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__6127\,
            I => \N__6120\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__6126\,
            I => \N__6117\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__6125\,
            I => \N__6113\
        );

    \I__1429\ : Span4Mux_h
    port map (
            O => \N__6120\,
            I => \N__6103\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6098\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6098\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6093\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6093\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6090\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6086\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6109\,
            I => \N__6083\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6108\,
            I => \N__6080\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6075\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6075\
        );

    \I__1418\ : Span4Mux_h
    port map (
            O => \N__6103\,
            I => \N__6070\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6098\,
            I => \N__6070\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6093\,
            I => \N__6067\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6064\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6089\,
            I => \N__6061\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6086\,
            I => \N__6058\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6055\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6080\,
            I => \N__6050\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6075\,
            I => \N__6050\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__6070\,
            I => \N__6041\
        );

    \I__1408\ : Span4Mux_v
    port map (
            O => \N__6067\,
            I => \N__6041\
        );

    \I__1407\ : Span4Mux_h
    port map (
            O => \N__6064\,
            I => \N__6041\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6041\
        );

    \I__1405\ : Span4Mux_v
    port map (
            O => \N__6058\,
            I => \N__6038\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__6055\,
            I => \N__6035\
        );

    \I__1403\ : Span4Mux_v
    port map (
            O => \N__6050\,
            I => \N__6032\
        );

    \I__1402\ : Span4Mux_v
    port map (
            O => \N__6041\,
            I => \N__6029\
        );

    \I__1401\ : Sp12to4
    port map (
            O => \N__6038\,
            I => \N__6026\
        );

    \I__1400\ : Span12Mux_v
    port map (
            O => \N__6035\,
            I => \N__6021\
        );

    \I__1399\ : Sp12to4
    port map (
            O => \N__6032\,
            I => \N__6021\
        );

    \I__1398\ : Sp12to4
    port map (
            O => \N__6029\,
            I => \N__6018\
        );

    \I__1397\ : Span12Mux_h
    port map (
            O => \N__6026\,
            I => \N__6015\
        );

    \I__1396\ : Span12Mux_v
    port map (
            O => \N__6021\,
            I => \N__6012\
        );

    \I__1395\ : Span12Mux_h
    port map (
            O => \N__6018\,
            I => \N__6009\
        );

    \I__1394\ : Span12Mux_v
    port map (
            O => \N__6015\,
            I => \N__6006\
        );

    \I__1393\ : Span12Mux_h
    port map (
            O => \N__6012\,
            I => \N__6001\
        );

    \I__1392\ : Span12Mux_v
    port map (
            O => \N__6009\,
            I => \N__6001\
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__6006\,
            I => \RESETn_c\
        );

    \I__1390\ : Odrv12
    port map (
            O => \N__6001\,
            I => \RESETn_c\
        );

    \I__1389\ : IoInMux
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__5993\,
            I => \N__5990\
        );

    \I__1387\ : Span4Mux_s3_v
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1386\ : Sp12to4
    port map (
            O => \N__5987\,
            I => \N__5984\
        );

    \I__1385\ : Span12Mux_h
    port map (
            O => \N__5984\,
            I => \N__5980\
        );

    \I__1384\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5977\
        );

    \I__1383\ : Span12Mux_v
    port map (
            O => \N__5980\,
            I => \N__5972\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__5977\,
            I => \N__5972\
        );

    \I__1381\ : Odrv12
    port map (
            O => \N__5972\,
            I => \nBUFEN_c\
        );

    \I__1380\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1378\ : Span4Mux_v
    port map (
            O => \N__5963\,
            I => \N__5960\
        );

    \I__1377\ : Sp12to4
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__1376\ : Span12Mux_h
    port map (
            O => \N__5957\,
            I => \N__5954\
        );

    \I__1375\ : Span12Mux_v
    port map (
            O => \N__5954\,
            I => \N__5951\
        );

    \I__1374\ : Odrv12
    port map (
            O => \N__5951\,
            I => \TACKn_in\
        );

    \I__1373\ : SRMux
    port map (
            O => \N__5948\,
            I => \N__5944\
        );

    \I__1372\ : SRMux
    port map (
            O => \N__5947\,
            I => \N__5940\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__5944\,
            I => \N__5937\
        );

    \I__1370\ : SRMux
    port map (
            O => \N__5943\,
            I => \N__5933\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5930\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__5937\,
            I => \N__5927\
        );

    \I__1367\ : SRMux
    port map (
            O => \N__5936\,
            I => \N__5924\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5921\
        );

    \I__1365\ : Span4Mux_v
    port map (
            O => \N__5930\,
            I => \N__5914\
        );

    \I__1364\ : Span4Mux_v
    port map (
            O => \N__5927\,
            I => \N__5914\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__5924\,
            I => \N__5914\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__5921\,
            I => \N__5911\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__5911\,
            I => \N__5903\
        );

    \I__1359\ : Span4Mux_h
    port map (
            O => \N__5908\,
            I => \N__5903\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__5903\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1357\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5894\
        );

    \I__1355\ : Span4Mux_v
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__5888\,
            I => \TACK_EN_i\
        );

    \I__1352\ : IoInMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1350\ : Span4Mux_s2_v
    port map (
            O => \N__5879\,
            I => \N__5876\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__5876\,
            I => \N__5873\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__5873\,
            I => \N__5870\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__5870\,
            I => \N_365_i\
        );

    \I__1346\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5856\
        );

    \I__1345\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5856\
        );

    \I__1344\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5849\
        );

    \I__1343\ : InMux
    port map (
            O => \N__5864\,
            I => \N__5849\
        );

    \I__1342\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5849\
        );

    \I__1341\ : InMux
    port map (
            O => \N__5862\,
            I => \N__5844\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5844\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5856\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5849\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__5844\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1336\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5834\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__5834\,
            I => \U409_CIA.CLKCIA6_0_a2_1\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__5831\,
            I => \N__5826\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__5830\,
            I => \N__5823\
        );

    \I__1332\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5819\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5826\,
            I => \N__5814\
        );

    \I__1330\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5814\
        );

    \I__1329\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5811\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__5819\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5814\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__5811\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5798\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5795\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5790\
        );

    \I__1322\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5790\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__5798\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__5795\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__5790\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1318\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5775\
        );

    \I__1317\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5775\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5772\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5780\,
            I => \N__5769\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5772\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5769\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5758\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5755\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5758\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5755\,
            I => \U409_CIA.CLKCIA8_0_a2_0\
        );

    \I__1307\ : SRMux
    port map (
            O => \N__5750\,
            I => \N__5746\
        );

    \I__1306\ : SRMux
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5737\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__1303\ : SRMux
    port map (
            O => \N__5742\,
            I => \N__5734\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__5737\,
            I => \N__5731\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__5734\,
            I => \N__5728\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__5731\,
            I => \RESETn_c_i\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__5728\,
            I => \RESETn_c_i\
        );

    \I__1298\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__5720\,
            I => \N__5717\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__5714\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5707\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__5698\,
            I => \N__5692\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__5695\,
            I => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__5692\,
            I => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__5687\,
            I => \N__5684\
        );

    \I__1285\ : InMux
    port map (
            O => \N__5684\,
            I => \N__5680\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5668\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5668\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5665\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5662\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5659\
        );

    \I__1278\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5655\
        );

    \I__1277\ : Span4Mux_h
    port map (
            O => \N__5668\,
            I => \N__5648\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5648\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5662\,
            I => \N__5648\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5645\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__5658\,
            I => \N__5641\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__5655\,
            I => \N__5638\
        );

    \I__1271\ : Span4Mux_v
    port map (
            O => \N__5648\,
            I => \N__5633\
        );

    \I__1270\ : Span4Mux_v
    port map (
            O => \N__5645\,
            I => \N__5633\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5630\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5627\
        );

    \I__1267\ : Span12Mux_h
    port map (
            O => \N__5638\,
            I => \N__5624\
        );

    \I__1266\ : Sp12to4
    port map (
            O => \N__5633\,
            I => \N__5621\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__5630\,
            I => \N__5616\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5627\,
            I => \N__5616\
        );

    \I__1263\ : Span12Mux_v
    port map (
            O => \N__5624\,
            I => \N__5613\
        );

    \I__1262\ : Span12Mux_h
    port map (
            O => \N__5621\,
            I => \N__5610\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__5616\,
            I => \N__5607\
        );

    \I__1260\ : Odrv12
    port map (
            O => \N__5613\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__5610\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__5607\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__5600\,
            I => \N__5597\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5594\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5594\,
            I => \N__5590\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5586\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__5590\,
            I => \N__5583\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5589\,
            I => \N__5580\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__5586\,
            I => \N__5577\
        );

    \I__1250\ : Span4Mux_v
    port map (
            O => \N__5583\,
            I => \N__5574\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5580\,
            I => \N__5571\
        );

    \I__1248\ : Span12Mux_h
    port map (
            O => \N__5577\,
            I => \N__5568\
        );

    \I__1247\ : Sp12to4
    port map (
            O => \N__5574\,
            I => \N__5563\
        );

    \I__1246\ : Span12Mux_v
    port map (
            O => \N__5571\,
            I => \N__5563\
        );

    \I__1245\ : Span12Mux_v
    port map (
            O => \N__5568\,
            I => \N__5558\
        );

    \I__1244\ : Span12Mux_h
    port map (
            O => \N__5563\,
            I => \N__5558\
        );

    \I__1243\ : Odrv12
    port map (
            O => \N__5558\,
            I => \OVL_c\
        );

    \I__1242\ : IoInMux
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__5552\,
            I => \N__5549\
        );

    \I__1240\ : Span4Mux_s3_v
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__1238\ : Sp12to4
    port map (
            O => \N__5543\,
            I => \N__5540\
        );

    \I__1237\ : Span12Mux_v
    port map (
            O => \N__5540\,
            I => \N__5536\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__1235\ : Odrv12
    port map (
            O => \N__5536\,
            I => \TACK_OUTn\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5533\,
            I => \TACK_OUTn\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5528\,
            I => \N__5524\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5527\,
            I => \N__5521\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__5524\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5521\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5513\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_0\
        );

    \I__1227\ : CascadeMux
    port map (
            O => \N__5510\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5507\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__5504\,
            I => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\
        );

    \I__1224\ : InMux
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5498\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5492\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1220\ : CascadeMux
    port map (
            O => \N__5489\,
            I => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\
        );

    \I__1219\ : CascadeMux
    port map (
            O => \N__5486\,
            I => \U409_CIA.N_20_cascade_\
        );

    \I__1218\ : CascadeMux
    port map (
            O => \N__5483\,
            I => \N__5473\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5470\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5481\,
            I => \N__5463\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5480\,
            I => \N__5463\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5463\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5454\
        );

    \I__1212\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5454\
        );

    \I__1211\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5454\
        );

    \I__1210\ : InMux
    port map (
            O => \N__5473\,
            I => \N__5454\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__5470\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5463\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5454\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__5447\,
            I => \U409_CIA.CLKCIAZ0_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5436\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5429\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5442\,
            I => \N__5429\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5441\,
            I => \N__5429\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5424\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5424\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5429\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5424\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1194\ : Span12Mux_s6_v
    port map (
            O => \N__5411\,
            I => \N__5407\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5410\,
            I => \N__5404\
        );

    \I__1192\ : Span12Mux_v
    port map (
            O => \N__5407\,
            I => \N__5400\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5404\,
            I => \N__5397\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5394\
        );

    \I__1189\ : Odrv12
    port map (
            O => \N__5400\,
            I => \CLKCIA_c\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__5397\,
            I => \CLKCIA_c\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5394\,
            I => \CLKCIA_c\
        );

    \I__1186\ : ClkMux
    port map (
            O => \N__5387\,
            I => \N__5375\
        );

    \I__1185\ : ClkMux
    port map (
            O => \N__5386\,
            I => \N__5375\
        );

    \I__1184\ : ClkMux
    port map (
            O => \N__5385\,
            I => \N__5375\
        );

    \I__1183\ : ClkMux
    port map (
            O => \N__5384\,
            I => \N__5375\
        );

    \I__1182\ : GlobalMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__1181\ : gio2CtrlBuf
    port map (
            O => \N__5372\,
            I => \CLK28_IN_c_g\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__5369\,
            I => \N__5365\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5357\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5362\,
            I => \N__5357\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__5357\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5351\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5337\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5337\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5346\,
            I => \N__5337\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5345\,
            I => \N__5332\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5332\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5337\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__5332\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5327\,
            I => \N__5316\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5316\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5316\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5311\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5311\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5316\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5311\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__5306\,
            I => \N__5301\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5305\,
            I => \N__5297\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5289\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5289\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5289\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5284\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5296\,
            I => \N__5284\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5289\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5284\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__5276\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5270\,
            I => \N__5261\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5256\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5256\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5253\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5246\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5246\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5246\
        );

    \I__1140\ : Odrv4
    port map (
            O => \N__5261\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5256\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5253\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5246\,
            I => \U409_TICK.TICK603_14\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5228\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5225\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5218\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5218\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5218\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5232\,
            I => \N__5213\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5231\,
            I => \N__5213\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5228\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5225\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5218\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5213\,
            I => \U409_TICK.TICK603_10\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__5204\,
            I => \N__5199\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__5203\,
            I => \N__5196\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5202\,
            I => \N__5189\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5199\,
            I => \N__5186\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5196\,
            I => \N__5183\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5195\,
            I => \N__5180\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5194\,
            I => \N__5175\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5193\,
            I => \N__5175\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5192\,
            I => \N__5170\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5170\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5186\,
            I => \N__5167\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__5183\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5180\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5175\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__5170\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1110\ : Odrv4
    port map (
            O => \N__5167\,
            I => \U409_TICK.TICK603_9\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5153\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5150\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__5150\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5147\,
            I => \N__5143\
        );

    \I__1105\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5140\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5137\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__1102\ : Odrv4
    port map (
            O => \N__5137\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__5134\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__1100\ : ClkMux
    port map (
            O => \N__5129\,
            I => \N__5093\
        );

    \I__1099\ : ClkMux
    port map (
            O => \N__5128\,
            I => \N__5093\
        );

    \I__1098\ : ClkMux
    port map (
            O => \N__5127\,
            I => \N__5093\
        );

    \I__1097\ : ClkMux
    port map (
            O => \N__5126\,
            I => \N__5093\
        );

    \I__1096\ : ClkMux
    port map (
            O => \N__5125\,
            I => \N__5093\
        );

    \I__1095\ : ClkMux
    port map (
            O => \N__5124\,
            I => \N__5093\
        );

    \I__1094\ : ClkMux
    port map (
            O => \N__5123\,
            I => \N__5093\
        );

    \I__1093\ : ClkMux
    port map (
            O => \N__5122\,
            I => \N__5093\
        );

    \I__1092\ : ClkMux
    port map (
            O => \N__5121\,
            I => \N__5093\
        );

    \I__1091\ : ClkMux
    port map (
            O => \N__5120\,
            I => \N__5093\
        );

    \I__1090\ : ClkMux
    port map (
            O => \N__5119\,
            I => \N__5093\
        );

    \I__1089\ : ClkMux
    port map (
            O => \N__5118\,
            I => \N__5093\
        );

    \I__1088\ : GlobalMux
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__1087\ : gio2CtrlBuf
    port map (
            O => \N__5090\,
            I => \CLK6_c_g\
        );

    \I__1086\ : InMux
    port map (
            O => \N__5087\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5084\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5081\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5075\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__5075\,
            I => \N__5072\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__5072\,
            I => \N__5067\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5062\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5070\,
            I => \N__5062\
        );

    \I__1078\ : Sp12to4
    port map (
            O => \N__5067\,
            I => \N__5057\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5062\,
            I => \N__5057\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__5057\,
            I => \U409_CIA.g0Z0Z_14\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__5054\,
            I => \N__5050\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5045\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5040\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5049\,
            I => \N__5040\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5048\,
            I => \N__5037\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5045\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5040\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5037\,
            I => \U409_CIA.VMAZ0\
        );

    \I__1067\ : CascadeMux
    port map (
            O => \N__5030\,
            I => \N__5026\
        );

    \I__1066\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5020\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5026\,
            I => \N__5020\
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__5025\,
            I => \N__5017\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5020\,
            I => \N__5014\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5011\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__5014\,
            I => \N__5006\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__5011\,
            I => \N__5006\
        );

    \I__1059\ : Span4Mux_v
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__1058\ : Sp12to4
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__1057\ : Span12Mux_h
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__4997\,
            I => \U409_CIA.g0Z0Z_13\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__4991\,
            I => \N__4986\
        );

    \I__1053\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4981\
        );

    \I__1052\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4981\
        );

    \I__1051\ : Odrv4
    port map (
            O => \N__4986\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__4981\,
            I => \U409_CIA.CIA_HOLDZ0\
        );

    \I__1049\ : CascadeMux
    port map (
            O => \N__4976\,
            I => \N__4970\
        );

    \I__1048\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4967\
        );

    \I__1047\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4960\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4960\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4970\,
            I => \N__4960\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__4967\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__4960\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4948\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4954\,
            I => \N__4939\
        );

    \I__1040\ : InMux
    port map (
            O => \N__4953\,
            I => \N__4939\
        );

    \I__1039\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4939\
        );

    \I__1038\ : InMux
    port map (
            O => \N__4951\,
            I => \N__4939\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4948\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__4928\,
            I => \U409_TRANSFER_ACK.N_105\
        );

    \I__1032\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4919\
        );

    \I__1031\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4912\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4912\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4922\,
            I => \N__4912\
        );

    \I__1028\ : LocalMux
    port map (
            O => \N__4919\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__4912\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__1026\ : CascadeMux
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4895\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4903\,
            I => \N__4895\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4902\,
            I => \N__4895\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__4895\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__1021\ : InMux
    port map (
            O => \N__4892\,
            I => \N__4887\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4882\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4882\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__4887\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__4882\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__1016\ : InMux
    port map (
            O => \N__4877\,
            I => \N__4871\
        );

    \I__1015\ : InMux
    port map (
            O => \N__4876\,
            I => \N__4871\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4871\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__1013\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4864\
        );

    \I__1012\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4861\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4861\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__4858\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4849\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4846\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__4849\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1005\ : LocalMux
    port map (
            O => \N__4846\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4837\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4834\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4837\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__4834\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1000\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4825\
        );

    \I__999\ : InMux
    port map (
            O => \N__4828\,
            I => \N__4822\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__4825\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__4822\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__995\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4811\,
            I => \N__4807\
        );

    \I__993\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4804\
        );

    \I__992\ : Odrv4
    port map (
            O => \N__4807\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4804\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__4799\,
            I => \N__4795\
        );

    \I__989\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4792\
        );

    \I__988\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4789\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4792\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__4789\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__4784\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__984\ : InMux
    port map (
            O => \N__4781\,
            I => \N__4778\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__4778\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__982\ : InMux
    port map (
            O => \N__4775\,
            I => \N__4771\
        );

    \I__981\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4768\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__4771\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__4768\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__978\ : InMux
    port map (
            O => \N__4763\,
            I => \N__4759\
        );

    \I__977\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4759\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__4756\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__974\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4747\
        );

    \I__973\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4744\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4747\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4744\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4739\,
            I => \N__4733\
        );

    \I__969\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4730\
        );

    \I__968\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4725\
        );

    \I__967\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4725\
        );

    \I__966\ : InMux
    port map (
            O => \N__4733\,
            I => \N__4722\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4730\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4725\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4722\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__962\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4712\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__4712\,
            I => \U409_TICK.TICK603_11\
        );

    \I__960\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4705\
        );

    \I__959\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4705\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4702\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__4697\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__955\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4690\
        );

    \I__954\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4690\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4687\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__4682\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__950\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4676\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4676\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__948\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4669\
        );

    \I__947\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4666\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4669\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4666\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__944\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4655\
        );

    \I__943\ : InMux
    port map (
            O => \N__4660\,
            I => \N__4655\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4652\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4652\,
            I => \CIA_ENABLEm\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__4649\,
            I => \U409_CIA.N_9_cascade_\
        );

    \I__939\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4643\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4643\,
            I => \N__4640\
        );

    \I__937\ : Span4Mux_v
    port map (
            O => \N__4640\,
            I => \N__4637\
        );

    \I__936\ : Sp12to4
    port map (
            O => \N__4637\,
            I => \N__4634\
        );

    \I__935\ : Span12Mux_h
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__934\ : Odrv12
    port map (
            O => \N__4631\,
            I => \A_c_13\
        );

    \I__933\ : IoInMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4625\,
            I => \N__4622\
        );

    \I__931\ : Span12Mux_s4_h
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__930\ : Span12Mux_h
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__929\ : Odrv12
    port map (
            O => \N__4616\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS1_i\
        );

    \I__928\ : IoInMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__926\ : Span12Mux_s4_v
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__925\ : Odrv12
    port map (
            O => \N__4604\,
            I => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\
        );

    \I__924\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__4598\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__922\ : IoInMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__920\ : Span4Mux_s3_v
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__919\ : Sp12to4
    port map (
            O => \N__4586\,
            I => \N__4583\
        );

    \I__918\ : Span12Mux_h
    port map (
            O => \N__4583\,
            I => \N__4579\
        );

    \I__917\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4576\
        );

    \I__916\ : Odrv12
    port map (
            O => \N__4579\,
            I => \TICK60_c\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__4576\,
            I => \TICK60_c\
        );

    \I__914\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4567\
        );

    \I__913\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4567\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__4564\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__910\ : InMux
    port map (
            O => \N__4559\,
            I => \N__4555\
        );

    \I__909\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4552\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4555\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__4552\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__4547\,
            I => \N__4543\
        );

    \I__905\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4537\
        );

    \I__904\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4537\
        );

    \I__903\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4534\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4537\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4534\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__900\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4525\
        );

    \I__899\ : InMux
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4525\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4522\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__895\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__4511\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__892\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4501\
        );

    \I__891\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4498\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4501\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__4498\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__888\ : CascadeMux
    port map (
            O => \N__4493\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__4490\,
            I => \U409_TRANSFER_ACK.N_105_cascade_\
        );

    \I__886\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4484\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4484\,
            I => \U409_TRANSFER_ACK.m9_bm\
        );

    \I__884\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4475\
        );

    \I__883\ : InMux
    port map (
            O => \N__4480\,
            I => \N__4475\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4475\,
            I => \U409_TRANSFER_ACK.N_4\
        );

    \I__881\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4469\,
            I => \N__4465\
        );

    \I__879\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4461\
        );

    \I__878\ : Span4Mux_v
    port map (
            O => \N__4465\,
            I => \N__4454\
        );

    \I__877\ : InMux
    port map (
            O => \N__4464\,
            I => \N__4451\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4461\,
            I => \N__4448\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4460\,
            I => \N__4445\
        );

    \I__874\ : InMux
    port map (
            O => \N__4459\,
            I => \N__4442\
        );

    \I__873\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4439\
        );

    \I__872\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4436\
        );

    \I__871\ : Sp12to4
    port map (
            O => \N__4454\,
            I => \N__4431\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4431\
        );

    \I__869\ : Span4Mux_v
    port map (
            O => \N__4448\,
            I => \N__4428\
        );

    \I__868\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4425\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4420\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4439\,
            I => \N__4420\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4436\,
            I => \N__4417\
        );

    \I__864\ : Span12Mux_h
    port map (
            O => \N__4431\,
            I => \N__4412\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__4428\,
            I => \N__4412\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4425\,
            I => \N__4405\
        );

    \I__861\ : Sp12to4
    port map (
            O => \N__4420\,
            I => \N__4405\
        );

    \I__860\ : Sp12to4
    port map (
            O => \N__4417\,
            I => \N__4405\
        );

    \I__859\ : Span12Mux_v
    port map (
            O => \N__4412\,
            I => \N__4402\
        );

    \I__858\ : Span12Mux_v
    port map (
            O => \N__4405\,
            I => \N__4399\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__4402\,
            I => \A_c_22\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__4399\,
            I => \A_c_22\
        );

    \I__855\ : InMux
    port map (
            O => \N__4394\,
            I => \N__4389\
        );

    \I__854\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4386\
        );

    \I__853\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4381\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__4389\,
            I => \N__4378\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4386\,
            I => \N__4375\
        );

    \I__850\ : InMux
    port map (
            O => \N__4385\,
            I => \N__4372\
        );

    \I__849\ : InMux
    port map (
            O => \N__4384\,
            I => \N__4368\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4381\,
            I => \N__4362\
        );

    \I__847\ : Span4Mux_v
    port map (
            O => \N__4378\,
            I => \N__4355\
        );

    \I__846\ : Span4Mux_h
    port map (
            O => \N__4375\,
            I => \N__4355\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4372\,
            I => \N__4355\
        );

    \I__844\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4352\
        );

    \I__843\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4349\
        );

    \I__842\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4346\
        );

    \I__841\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4343\
        );

    \I__840\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4340\
        );

    \I__839\ : Span4Mux_v
    port map (
            O => \N__4362\,
            I => \N__4335\
        );

    \I__838\ : Span4Mux_v
    port map (
            O => \N__4355\,
            I => \N__4335\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4352\,
            I => \N__4332\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__4349\,
            I => \N__4329\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4346\,
            I => \N__4326\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4321\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4340\,
            I => \N__4321\
        );

    \I__832\ : Span4Mux_h
    port map (
            O => \N__4335\,
            I => \N__4316\
        );

    \I__831\ : Span4Mux_v
    port map (
            O => \N__4332\,
            I => \N__4316\
        );

    \I__830\ : Span4Mux_v
    port map (
            O => \N__4329\,
            I => \N__4309\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__4326\,
            I => \N__4309\
        );

    \I__828\ : Span4Mux_v
    port map (
            O => \N__4321\,
            I => \N__4309\
        );

    \I__827\ : Sp12to4
    port map (
            O => \N__4316\,
            I => \N__4304\
        );

    \I__826\ : Sp12to4
    port map (
            O => \N__4309\,
            I => \N__4304\
        );

    \I__825\ : Odrv12
    port map (
            O => \N__4304\,
            I => \A_c_23\
        );

    \I__824\ : InMux
    port map (
            O => \N__4301\,
            I => \N__4297\
        );

    \I__823\ : InMux
    port map (
            O => \N__4300\,
            I => \N__4293\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__4297\,
            I => \N__4289\
        );

    \I__821\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4286\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4293\,
            I => \N__4283\
        );

    \I__819\ : CascadeMux
    port map (
            O => \N__4292\,
            I => \N__4278\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__4289\,
            I => \N__4275\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4272\
        );

    \I__816\ : Span4Mux_h
    port map (
            O => \N__4283\,
            I => \N__4269\
        );

    \I__815\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4266\
        );

    \I__814\ : InMux
    port map (
            O => \N__4281\,
            I => \N__4261\
        );

    \I__813\ : InMux
    port map (
            O => \N__4278\,
            I => \N__4261\
        );

    \I__812\ : Span4Mux_v
    port map (
            O => \N__4275\,
            I => \N__4258\
        );

    \I__811\ : Span4Mux_v
    port map (
            O => \N__4272\,
            I => \N__4255\
        );

    \I__810\ : Span4Mux_h
    port map (
            O => \N__4269\,
            I => \N__4248\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4266\,
            I => \N__4248\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4261\,
            I => \N__4248\
        );

    \I__807\ : Span4Mux_h
    port map (
            O => \N__4258\,
            I => \N__4245\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__4255\,
            I => \N__4240\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__4248\,
            I => \N__4240\
        );

    \I__804\ : Sp12to4
    port map (
            O => \N__4245\,
            I => \N__4235\
        );

    \I__803\ : Sp12to4
    port map (
            O => \N__4240\,
            I => \N__4235\
        );

    \I__802\ : Odrv12
    port map (
            O => \N__4235\,
            I => \A_c_21\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__800\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4225\
        );

    \I__799\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4222\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N__4217\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4222\,
            I => \N__4217\
        );

    \I__796\ : Odrv12
    port map (
            O => \N__4217\,
            I => \U409_ADDRESS_DECODE.LOWROMZ0\
        );

    \I__795\ : CascadeMux
    port map (
            O => \N__4214\,
            I => \N__4210\
        );

    \I__794\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__793\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4204\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4201\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N__4198\
        );

    \I__790\ : Span12Mux_v
    port map (
            O => \N__4201\,
            I => \N__4195\
        );

    \I__789\ : Span4Mux_h
    port map (
            O => \N__4198\,
            I => \N__4192\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__4195\,
            I => \U409_ADDRESS_DECODE.HIROMZ0\
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4192\,
            I => \U409_ADDRESS_DECODE.HIROMZ0\
        );

    \I__786\ : IoInMux
    port map (
            O => \N__4187\,
            I => \N__4184\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4184\,
            I => \N__4181\
        );

    \I__784\ : Span4Mux_s0_v
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__783\ : Span4Mux_v
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__782\ : Sp12to4
    port map (
            O => \N__4175\,
            I => \N__4172\
        );

    \I__781\ : Span12Mux_h
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__780\ : Odrv12
    port map (
            O => \N__4169\,
            I => \ROMENm_i\
        );

    \I__779\ : InMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__777\ : Span4Mux_v
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__775\ : Odrv4
    port map (
            O => \N__4154\,
            I => \AUTOVECTORm\
        );

    \I__774\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4145\
        );

    \I__773\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4145\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__4145\,
            I => \N__4142\
        );

    \I__771\ : Span4Mux_v
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__4139\,
            I => \N__4135\
        );

    \I__769\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4132\
        );

    \I__768\ : Sp12to4
    port map (
            O => \N__4135\,
            I => \N__4127\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4127\
        );

    \I__766\ : Span12Mux_h
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__765\ : Span12Mux_v
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__4121\,
            I => \TSn_c\
        );

    \I__763\ : IoInMux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4111\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__4114\,
            I => \N__4107\
        );

    \I__760\ : IoSpan4Mux
    port map (
            O => \N__4111\,
            I => \N__4102\
        );

    \I__759\ : InMux
    port map (
            O => \N__4110\,
            I => \N__4099\
        );

    \I__758\ : InMux
    port map (
            O => \N__4107\,
            I => \N__4096\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__4106\,
            I => \N__4093\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__4105\,
            I => \N__4090\
        );

    \I__755\ : Span4Mux_s0_v
    port map (
            O => \N__4102\,
            I => \N__4087\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4099\,
            I => \N__4084\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4096\,
            I => \N__4081\
        );

    \I__752\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4078\
        );

    \I__751\ : InMux
    port map (
            O => \N__4090\,
            I => \N__4075\
        );

    \I__750\ : Sp12to4
    port map (
            O => \N__4087\,
            I => \N__4072\
        );

    \I__749\ : Span4Mux_v
    port map (
            O => \N__4084\,
            I => \N__4065\
        );

    \I__748\ : Span4Mux_v
    port map (
            O => \N__4081\,
            I => \N__4065\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4078\,
            I => \N__4065\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4075\,
            I => \N__4062\
        );

    \I__745\ : Span12Mux_v
    port map (
            O => \N__4072\,
            I => \N__4055\
        );

    \I__744\ : Sp12to4
    port map (
            O => \N__4065\,
            I => \N__4055\
        );

    \I__743\ : Sp12to4
    port map (
            O => \N__4062\,
            I => \N__4055\
        );

    \I__742\ : Span12Mux_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__741\ : Odrv12
    port map (
            O => \N__4052\,
            I => \CLK40_IN_c\
        );

    \I__740\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__738\ : Odrv4
    port map (
            O => \N__4043\,
            I => \ROMENm\
        );

    \I__737\ : IoInMux
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__735\ : Span4Mux_s3_v
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__734\ : Span4Mux_h
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__4028\,
            I => \CONSTANT_ONE_NET\
        );

    \I__732\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__730\ : Span12Mux_s10_v
    port map (
            O => \N__4019\,
            I => \N__4016\
        );

    \I__729\ : Span12Mux_h
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__728\ : Odrv12
    port map (
            O => \N__4013\,
            I => \A_c_12\
        );

    \I__727\ : IoInMux
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4007\,
            I => \N__4004\
        );

    \I__725\ : IoSpan4Mux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__724\ : Span4Mux_s3_h
    port map (
            O => \N__4001\,
            I => \N__3998\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__722\ : Span4Mux_h
    port map (
            O => \N__3995\,
            I => \N__3992\
        );

    \I__721\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__720\ : Odrv12
    port map (
            O => \N__3989\,
            I => \U409_ADDRESS_DECODE_un1_nCIACS0_i\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__3986\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__3983\,
            I => \N__3979\
        );

    \I__717\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3976\
        );

    \I__716\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3973\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__3976\,
            I => \N__3965\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__3973\,
            I => \N__3962\
        );

    \I__713\ : InMux
    port map (
            O => \N__3972\,
            I => \N__3951\
        );

    \I__712\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3951\
        );

    \I__711\ : InMux
    port map (
            O => \N__3970\,
            I => \N__3951\
        );

    \I__710\ : InMux
    port map (
            O => \N__3969\,
            I => \N__3951\
        );

    \I__709\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3951\
        );

    \I__708\ : Odrv4
    port map (
            O => \N__3965\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__707\ : Odrv4
    port map (
            O => \N__3962\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__3951\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__705\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3937\
        );

    \I__704\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3934\
        );

    \I__703\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3927\
        );

    \I__702\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3927\
        );

    \I__701\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3927\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3937\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__3934\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3927\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__697\ : InMux
    port map (
            O => \N__3920\,
            I => \N__3914\
        );

    \I__696\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3911\
        );

    \I__695\ : InMux
    port map (
            O => \N__3918\,
            I => \N__3906\
        );

    \I__694\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3906\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__3914\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3911\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__3906\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__690\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3896\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\
        );

    \I__688\ : InMux
    port map (
            O => \N__3893\,
            I => \N__3888\
        );

    \I__687\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3883\
        );

    \I__686\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3883\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__3888\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__3883\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__3878\,
            I => \U409_TRANSFER_ACK.m9_am_cascade_\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__3875\,
            I => \U409_TRANSFER_ACK.i6_mux_0_cascade_\
        );

    \I__681\ : CascadeMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__680\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3866\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__678\ : InMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__3857\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\
        );

    \I__675\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3851\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3\
        );

    \I__673\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3844\
        );

    \I__672\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3840\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__3844\,
            I => \N__3837\
        );

    \I__670\ : InMux
    port map (
            O => \N__3843\,
            I => \N__3834\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3840\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__668\ : Odrv4
    port map (
            O => \N__3837\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3834\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__666\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3821\
        );

    \I__665\ : InMux
    port map (
            O => \N__3826\,
            I => \N__3818\
        );

    \I__664\ : InMux
    port map (
            O => \N__3825\,
            I => \N__3815\
        );

    \I__663\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3812\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__3821\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__3818\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3815\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3812\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__658\ : CascadeMux
    port map (
            O => \N__3803\,
            I => \N__3798\
        );

    \I__657\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3792\
        );

    \I__656\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3792\
        );

    \I__655\ : InMux
    port map (
            O => \N__3798\,
            I => \N__3787\
        );

    \I__654\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3787\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3792\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3787\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__3782\,
            I => \N__3777\
        );

    \I__650\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3773\
        );

    \I__649\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3770\
        );

    \I__648\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3767\
        );

    \I__647\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3764\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__3773\,
            I => \N__3761\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3756\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__3767\,
            I => \N__3756\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3764\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__3761\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__3756\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__640\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3742\
        );

    \I__639\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3737\
        );

    \I__638\ : InMux
    port map (
            O => \N__3747\,
            I => \N__3737\
        );

    \I__637\ : InMux
    port map (
            O => \N__3746\,
            I => \N__3734\
        );

    \I__636\ : InMux
    port map (
            O => \N__3745\,
            I => \N__3731\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3742\,
            I => \N__3728\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3737\,
            I => \N__3723\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3734\,
            I => \N__3723\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__3731\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__3728\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__3723\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__3716\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__627\ : InMux
    port map (
            O => \N__3710\,
            I => \N__3704\
        );

    \I__626\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3704\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3704\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__3701\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__3698\,
            I => \N__3694\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3697\,
            I => \N__3689\
        );

    \I__621\ : InMux
    port map (
            O => \N__3694\,
            I => \N__3683\
        );

    \I__620\ : InMux
    port map (
            O => \N__3693\,
            I => \N__3683\
        );

    \I__619\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3676\
        );

    \I__618\ : InMux
    port map (
            O => \N__3689\,
            I => \N__3676\
        );

    \I__617\ : InMux
    port map (
            O => \N__3688\,
            I => \N__3676\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__3683\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3676\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__614\ : InMux
    port map (
            O => \N__3671\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__613\ : InMux
    port map (
            O => \N__3668\,
            I => \bfn_11_6_0_\
        );

    \I__612\ : InMux
    port map (
            O => \N__3665\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__611\ : InMux
    port map (
            O => \N__3662\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__610\ : InMux
    port map (
            O => \N__3659\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__609\ : InMux
    port map (
            O => \N__3656\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__608\ : InMux
    port map (
            O => \N__3653\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__607\ : InMux
    port map (
            O => \N__3650\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__606\ : InMux
    port map (
            O => \N__3647\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__605\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__3638\,
            I => \N__3633\
        );

    \I__602\ : InMux
    port map (
            O => \N__3637\,
            I => \N__3630\
        );

    \I__601\ : InMux
    port map (
            O => \N__3636\,
            I => \N__3627\
        );

    \I__600\ : Span4Mux_h
    port map (
            O => \N__3633\,
            I => \N__3624\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3630\,
            I => \N__3621\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3627\,
            I => \N__3618\
        );

    \I__597\ : Odrv4
    port map (
            O => \N__3624\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__596\ : Odrv12
    port map (
            O => \N__3621\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__595\ : Odrv12
    port map (
            O => \N__3618\,
            I => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\
        );

    \I__594\ : IoInMux
    port map (
            O => \N__3611\,
            I => \N__3608\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3608\,
            I => \N__3605\
        );

    \I__592\ : IoSpan4Mux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__591\ : Sp12to4
    port map (
            O => \N__3602\,
            I => \N__3599\
        );

    \I__590\ : Span12Mux_s6_v
    port map (
            O => \N__3599\,
            I => \N__3596\
        );

    \I__589\ : Span12Mux_h
    port map (
            O => \N__3596\,
            I => \N__3593\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__3593\,
            I => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\
        );

    \I__587\ : InMux
    port map (
            O => \N__3590\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__586\ : InMux
    port map (
            O => \N__3587\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__585\ : InMux
    port map (
            O => \N__3584\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__584\ : InMux
    port map (
            O => \N__3581\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__583\ : InMux
    port map (
            O => \N__3578\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__582\ : InMux
    port map (
            O => \N__3575\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__581\ : IoInMux
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__579\ : Span4Mux_s1_v
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__578\ : Sp12to4
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__577\ : Span12Mux_h
    port map (
            O => \N__3560\,
            I => \N__3556\
        );

    \I__576\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3553\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__3556\,
            I => \TICK50_c\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__3553\,
            I => \TICK50_c\
        );

    \I__573\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3533\
        );

    \I__572\ : InMux
    port map (
            O => \N__3547\,
            I => \N__3533\
        );

    \I__571\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3533\
        );

    \I__570\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3533\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__3544\,
            I => \N__3530\
        );

    \I__568\ : InMux
    port map (
            O => \N__3543\,
            I => \N__3526\
        );

    \I__567\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3523\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3533\,
            I => \N__3520\
        );

    \I__565\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3515\
        );

    \I__564\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3515\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3526\,
            I => \U409_TICK.TICK503_14\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3523\,
            I => \U409_TICK.TICK503_14\
        );

    \I__561\ : Odrv4
    port map (
            O => \N__3520\,
            I => \U409_TICK.TICK503_14\
        );

    \I__560\ : LocalMux
    port map (
            O => \N__3515\,
            I => \U409_TICK.TICK503_14\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3506\,
            I => \N__3503\
        );

    \I__558\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3493\
        );

    \I__557\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3486\
        );

    \I__556\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3486\
        );

    \I__555\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3486\
        );

    \I__554\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3483\
        );

    \I__553\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3476\
        );

    \I__552\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3476\
        );

    \I__551\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3476\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3493\,
            I => \U409_TICK.TICK503_9\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3486\,
            I => \U409_TICK.TICK503_9\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3483\,
            I => \U409_TICK.TICK503_9\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__3476\,
            I => \U409_TICK.TICK503_9\
        );

    \I__546\ : CascadeMux
    port map (
            O => \N__3467\,
            I => \N__3461\
        );

    \I__545\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \N__3457\
        );

    \I__544\ : CascadeMux
    port map (
            O => \N__3465\,
            I => \N__3454\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3464\,
            I => \N__3451\
        );

    \I__542\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3445\
        );

    \I__541\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3442\
        );

    \I__540\ : InMux
    port map (
            O => \N__3457\,
            I => \N__3435\
        );

    \I__539\ : InMux
    port map (
            O => \N__3454\,
            I => \N__3435\
        );

    \I__538\ : InMux
    port map (
            O => \N__3451\,
            I => \N__3435\
        );

    \I__537\ : InMux
    port map (
            O => \N__3450\,
            I => \N__3432\
        );

    \I__536\ : InMux
    port map (
            O => \N__3449\,
            I => \N__3427\
        );

    \I__535\ : InMux
    port map (
            O => \N__3448\,
            I => \N__3427\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3445\,
            I => \U409_TICK.TICK503_10\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3442\,
            I => \U409_TICK.TICK503_10\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3435\,
            I => \U409_TICK.TICK503_10\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3432\,
            I => \U409_TICK.TICK503_10\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3427\,
            I => \U409_TICK.TICK503_10\
        );

    \I__529\ : InMux
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3413\,
            I => \N__3410\
        );

    \I__527\ : Odrv4
    port map (
            O => \N__3410\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__526\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3403\
        );

    \I__525\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3400\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3403\,
            I => \N__3397\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3400\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3397\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__521\ : InMux
    port map (
            O => \N__3392\,
            I => \N__3386\
        );

    \I__520\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3386\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__3383\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__3380\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__515\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3368\
        );

    \I__514\ : InMux
    port map (
            O => \N__3373\,
            I => \N__3368\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3368\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__512\ : InMux
    port map (
            O => \N__3365\,
            I => \N__3362\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3362\,
            I => \U409_TICK.TICK503_11\
        );

    \I__510\ : InMux
    port map (
            O => \N__3359\,
            I => \N__3355\
        );

    \I__509\ : InMux
    port map (
            O => \N__3358\,
            I => \N__3352\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__3355\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__3352\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__3347\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__505\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3341\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3341\,
            I => \N__3337\
        );

    \I__503\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3334\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__3337\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__3334\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__3329\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__499\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3323\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3323\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3320\,
            I => \N__3316\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3319\,
            I => \N__3313\
        );

    \I__495\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3307\
        );

    \I__494\ : InMux
    port map (
            O => \N__3313\,
            I => \N__3307\
        );

    \I__493\ : InMux
    port map (
            O => \N__3312\,
            I => \N__3304\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3307\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3304\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3299\,
            I => \N__3293\
        );

    \I__489\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3286\
        );

    \I__488\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3286\
        );

    \I__487\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3286\
        );

    \I__486\ : InMux
    port map (
            O => \N__3293\,
            I => \N__3283\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3286\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3283\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__483\ : InMux
    port map (
            O => \N__3278\,
            I => \N__3275\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3275\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__481\ : CascadeMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__480\ : InMux
    port map (
            O => \N__3269\,
            I => \N__3265\
        );

    \I__479\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3262\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3265\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3262\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__3257\,
            I => \N__3254\
        );

    \I__475\ : InMux
    port map (
            O => \N__3254\,
            I => \N__3251\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3251\,
            I => \N__3247\
        );

    \I__473\ : InMux
    port map (
            O => \N__3250\,
            I => \N__3244\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__3247\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3244\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__3239\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__469\ : InMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3233\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__467\ : InMux
    port map (
            O => \N__3230\,
            I => \N__3226\
        );

    \I__466\ : InMux
    port map (
            O => \N__3229\,
            I => \N__3223\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3226\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__3223\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__463\ : InMux
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3215\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__461\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3208\
        );

    \I__460\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3205\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3208\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3205\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__457\ : InMux
    port map (
            O => \N__3200\,
            I => \N__3197\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3197\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__455\ : InMux
    port map (
            O => \N__3194\,
            I => \N__3190\
        );

    \I__454\ : InMux
    port map (
            O => \N__3193\,
            I => \N__3187\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3190\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3187\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__451\ : InMux
    port map (
            O => \N__3182\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__450\ : InMux
    port map (
            O => \N__3179\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__449\ : InMux
    port map (
            O => \N__3176\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__448\ : InMux
    port map (
            O => \N__3173\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__447\ : InMux
    port map (
            O => \N__3170\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__446\ : InMux
    port map (
            O => \N__3167\,
            I => \N__3163\
        );

    \I__445\ : InMux
    port map (
            O => \N__3166\,
            I => \N__3160\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3163\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3160\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__442\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3151\
        );

    \I__441\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3148\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3151\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3148\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__438\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3139\
        );

    \I__437\ : InMux
    port map (
            O => \N__3142\,
            I => \N__3136\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3139\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3136\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__434\ : InMux
    port map (
            O => \N__3131\,
            I => \N__3127\
        );

    \I__433\ : InMux
    port map (
            O => \N__3130\,
            I => \N__3124\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3127\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3124\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__430\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3115\
        );

    \I__429\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3112\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3115\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3112\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3107\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__425\ : InMux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3101\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__423\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3094\
        );

    \I__422\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3091\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3094\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3091\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__419\ : InMux
    port map (
            O => \N__3086\,
            I => \N__3082\
        );

    \I__418\ : InMux
    port map (
            O => \N__3085\,
            I => \N__3079\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3082\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3079\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__415\ : InMux
    port map (
            O => \N__3074\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__414\ : InMux
    port map (
            O => \N__3071\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__413\ : InMux
    port map (
            O => \N__3068\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__412\ : InMux
    port map (
            O => \N__3065\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__411\ : InMux
    port map (
            O => \N__3062\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__410\ : InMux
    port map (
            O => \N__3059\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__409\ : InMux
    port map (
            O => \N__3056\,
            I => \bfn_8_6_0_\
        );

    \I__408\ : InMux
    port map (
            O => \N__3053\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__407\ : InMux
    port map (
            O => \N__3050\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__405\ : InMux
    port map (
            O => \N__3044\,
            I => \N__3038\
        );

    \I__404\ : InMux
    port map (
            O => \N__3043\,
            I => \N__3038\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3038\,
            I => \N__3034\
        );

    \I__402\ : InMux
    port map (
            O => \N__3037\,
            I => \N__3031\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__3034\,
            I => \N__3026\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3031\,
            I => \N__3026\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__3023\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_6\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__396\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3014\,
            I => \N__3010\
        );

    \I__394\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3007\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__3010\,
            I => \N__3004\
        );

    \I__392\ : LocalMux
    port map (
            O => \N__3007\,
            I => \N__3001\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__3004\,
            I => \N__2994\
        );

    \I__390\ : Span4Mux_v
    port map (
            O => \N__3001\,
            I => \N__2994\
        );

    \I__389\ : InMux
    port map (
            O => \N__3000\,
            I => \N__2991\
        );

    \I__388\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2988\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__2994\,
            I => \N__2981\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2991\,
            I => \N__2981\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2988\,
            I => \N__2981\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__2981\,
            I => \A_c_20\
        );

    \I__383\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__381\ : Odrv12
    port map (
            O => \N__2972\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0\
        );

    \I__380\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2966\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__377\ : Span4Mux_v
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__376\ : IoSpan4Mux
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__375\ : Odrv4
    port map (
            O => \N__2954\,
            I => \TT_c_1\
        );

    \I__374\ : InMux
    port map (
            O => \N__2951\,
            I => \N__2948\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__372\ : Span4Mux_h
    port map (
            O => \N__2945\,
            I => \N__2942\
        );

    \I__371\ : Span4Mux_v
    port map (
            O => \N__2942\,
            I => \N__2939\
        );

    \I__370\ : Span4Mux_v
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__369\ : Odrv4
    port map (
            O => \N__2936\,
            I => \TT_c_0\
        );

    \I__368\ : InMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__2927\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\
        );

    \I__365\ : InMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__363\ : Span12Mux_v
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__362\ : Odrv12
    port map (
            O => \N__2915\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0\
        );

    \I__361\ : CascadeMux
    port map (
            O => \N__2912\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_cascade_\
        );

    \I__360\ : IoInMux
    port map (
            O => \N__2909\,
            I => \N__2906\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__358\ : Span12Mux_s9_v
    port map (
            O => \N__2903\,
            I => \N__2900\
        );

    \I__357\ : Odrv12
    port map (
            O => \N__2900\,
            I => \PORTSIZE_0_i\
        );

    \I__356\ : InMux
    port map (
            O => \N__2897\,
            I => \N__2894\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__2894\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_3\
        );

    \I__354\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2886\
        );

    \I__353\ : InMux
    port map (
            O => \N__2890\,
            I => \N__2883\
        );

    \I__352\ : InMux
    port map (
            O => \N__2889\,
            I => \N__2880\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__2886\,
            I => \N__2877\
        );

    \I__350\ : LocalMux
    port map (
            O => \N__2883\,
            I => \N__2872\
        );

    \I__349\ : LocalMux
    port map (
            O => \N__2880\,
            I => \N__2872\
        );

    \I__348\ : Span12Mux_h
    port map (
            O => \N__2877\,
            I => \N__2869\
        );

    \I__347\ : Span12Mux_h
    port map (
            O => \N__2872\,
            I => \N__2866\
        );

    \I__346\ : Span12Mux_v
    port map (
            O => \N__2869\,
            I => \N__2863\
        );

    \I__345\ : Span12Mux_v
    port map (
            O => \N__2866\,
            I => \N__2860\
        );

    \I__344\ : Odrv12
    port map (
            O => \N__2863\,
            I => \A_c_19\
        );

    \I__343\ : Odrv12
    port map (
            O => \N__2860\,
            I => \A_c_19\
        );

    \I__342\ : InMux
    port map (
            O => \N__2855\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2852\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2846\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__338\ : Span4Mux_v
    port map (
            O => \N__2843\,
            I => \N__2838\
        );

    \I__337\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2833\
        );

    \I__336\ : InMux
    port map (
            O => \N__2841\,
            I => \N__2833\
        );

    \I__335\ : Span4Mux_v
    port map (
            O => \N__2838\,
            I => \N__2828\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2833\,
            I => \N__2828\
        );

    \I__333\ : Span4Mux_v
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__332\ : Span4Mux_v
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__331\ : Span4Mux_h
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__330\ : Odrv4
    port map (
            O => \N__2819\,
            I => \A_c_26\
        );

    \I__329\ : InMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__2810\,
            I => \N__2805\
        );

    \I__326\ : InMux
    port map (
            O => \N__2809\,
            I => \N__2800\
        );

    \I__325\ : InMux
    port map (
            O => \N__2808\,
            I => \N__2800\
        );

    \I__324\ : Sp12to4
    port map (
            O => \N__2805\,
            I => \N__2795\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2800\,
            I => \N__2795\
        );

    \I__322\ : Odrv12
    port map (
            O => \N__2795\,
            I => \A_c_27\
        );

    \I__321\ : InMux
    port map (
            O => \N__2792\,
            I => \N__2789\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2789\,
            I => \N__2785\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2788\,
            I => \N__2781\
        );

    \I__318\ : Span4Mux_v
    port map (
            O => \N__2785\,
            I => \N__2778\
        );

    \I__317\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2773\
        );

    \I__316\ : InMux
    port map (
            O => \N__2781\,
            I => \N__2773\
        );

    \I__315\ : Sp12to4
    port map (
            O => \N__2778\,
            I => \N__2768\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2773\,
            I => \N__2768\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__2768\,
            I => \A_c_25\
        );

    \I__312\ : InMux
    port map (
            O => \N__2765\,
            I => \N__2760\
        );

    \I__311\ : InMux
    port map (
            O => \N__2764\,
            I => \N__2755\
        );

    \I__310\ : InMux
    port map (
            O => \N__2763\,
            I => \N__2755\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2760\,
            I => \N__2750\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2755\,
            I => \N__2750\
        );

    \I__307\ : Span4Mux_v
    port map (
            O => \N__2750\,
            I => \N__2747\
        );

    \I__306\ : Span4Mux_v
    port map (
            O => \N__2747\,
            I => \N__2744\
        );

    \I__305\ : Sp12to4
    port map (
            O => \N__2744\,
            I => \N__2741\
        );

    \I__304\ : Odrv12
    port map (
            O => \N__2741\,
            I => \A_c_24\
        );

    \I__303\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2735\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2735\,
            I => \N__2732\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__2732\,
            I => \U409_CIA.g0Z0Z_10\
        );

    \I__300\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2720\
        );

    \I__299\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2720\
        );

    \I__298\ : InMux
    port map (
            O => \N__2727\,
            I => \N__2720\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__2720\,
            I => \N__2717\
        );

    \I__296\ : Span4Mux_v
    port map (
            O => \N__2717\,
            I => \N__2714\
        );

    \I__295\ : Sp12to4
    port map (
            O => \N__2714\,
            I => \N__2711\
        );

    \I__294\ : Odrv12
    port map (
            O => \N__2711\,
            I => \A_c_31\
        );

    \I__293\ : InMux
    port map (
            O => \N__2708\,
            I => \N__2699\
        );

    \I__292\ : InMux
    port map (
            O => \N__2707\,
            I => \N__2699\
        );

    \I__291\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2699\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2699\,
            I => \N__2696\
        );

    \I__289\ : Span4Mux_v
    port map (
            O => \N__2696\,
            I => \N__2693\
        );

    \I__288\ : Span4Mux_v
    port map (
            O => \N__2693\,
            I => \N__2690\
        );

    \I__287\ : Sp12to4
    port map (
            O => \N__2690\,
            I => \N__2687\
        );

    \I__286\ : Odrv12
    port map (
            O => \N__2687\,
            I => \A_c_28\
        );

    \I__285\ : InMux
    port map (
            O => \N__2684\,
            I => \N__2680\
        );

    \I__284\ : CascadeMux
    port map (
            O => \N__2683\,
            I => \N__2677\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2680\,
            I => \N__2673\
        );

    \I__282\ : InMux
    port map (
            O => \N__2677\,
            I => \N__2668\
        );

    \I__281\ : InMux
    port map (
            O => \N__2676\,
            I => \N__2668\
        );

    \I__280\ : Span4Mux_h
    port map (
            O => \N__2673\,
            I => \N__2663\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2668\,
            I => \N__2663\
        );

    \I__278\ : Span4Mux_v
    port map (
            O => \N__2663\,
            I => \N__2660\
        );

    \I__277\ : Span4Mux_h
    port map (
            O => \N__2660\,
            I => \N__2657\
        );

    \I__276\ : Odrv4
    port map (
            O => \N__2657\,
            I => \A_c_30\
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__2654\,
            I => \N__2650\
        );

    \I__274\ : CascadeMux
    port map (
            O => \N__2653\,
            I => \N__2646\
        );

    \I__273\ : InMux
    port map (
            O => \N__2650\,
            I => \N__2639\
        );

    \I__272\ : InMux
    port map (
            O => \N__2649\,
            I => \N__2639\
        );

    \I__271\ : InMux
    port map (
            O => \N__2646\,
            I => \N__2639\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2639\,
            I => \N__2636\
        );

    \I__269\ : Span4Mux_h
    port map (
            O => \N__2636\,
            I => \N__2633\
        );

    \I__268\ : Span4Mux_v
    port map (
            O => \N__2633\,
            I => \N__2630\
        );

    \I__267\ : Odrv4
    port map (
            O => \N__2630\,
            I => \A_c_29\
        );

    \I__266\ : InMux
    port map (
            O => \N__2627\,
            I => \N__2624\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2624\,
            I => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\
        );

    \I__264\ : InMux
    port map (
            O => \N__2621\,
            I => \N__2618\
        );

    \I__263\ : LocalMux
    port map (
            O => \N__2618\,
            I => \U409_CIA.g0Z0Z_8\
        );

    \I__262\ : CascadeMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__261\ : InMux
    port map (
            O => \N__2612\,
            I => \N__2609\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2609\,
            I => \N__2605\
        );

    \I__259\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2602\
        );

    \I__258\ : Span4Mux_h
    port map (
            O => \N__2605\,
            I => \N__2597\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2602\,
            I => \N__2597\
        );

    \I__256\ : Span4Mux_v
    port map (
            O => \N__2597\,
            I => \N__2594\
        );

    \I__255\ : Span4Mux_h
    port map (
            O => \N__2594\,
            I => \N__2591\
        );

    \I__254\ : Span4Mux_v
    port map (
            O => \N__2591\,
            I => \N__2588\
        );

    \I__253\ : Odrv4
    port map (
            O => \N__2588\,
            I => \A_c_16\
        );

    \I__252\ : InMux
    port map (
            O => \N__2585\,
            I => \N__2582\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2582\,
            I => \U409_CIA.g0Z0Z_11\
        );

    \I__250\ : InMux
    port map (
            O => \N__2579\,
            I => \N__2576\
        );

    \I__249\ : LocalMux
    port map (
            O => \N__2576\,
            I => \N__2573\
        );

    \I__248\ : Span4Mux_h
    port map (
            O => \N__2573\,
            I => \N__2570\
        );

    \I__247\ : Odrv4
    port map (
            O => \N__2570\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\
        );

    \I__246\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2564\,
            I => \N__2561\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2561\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\
        );

    \I__243\ : CascadeMux
    port map (
            O => \N__2558\,
            I => \U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_\
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__2555\,
            I => \N__2551\
        );

    \I__241\ : InMux
    port map (
            O => \N__2554\,
            I => \N__2548\
        );

    \I__240\ : InMux
    port map (
            O => \N__2551\,
            I => \N__2545\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__2548\,
            I => \N__2540\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__2545\,
            I => \N__2540\
        );

    \I__237\ : Span4Mux_v
    port map (
            O => \N__2540\,
            I => \N__2537\
        );

    \I__236\ : Span4Mux_h
    port map (
            O => \N__2537\,
            I => \N__2534\
        );

    \I__235\ : Span4Mux_v
    port map (
            O => \N__2534\,
            I => \N__2531\
        );

    \I__234\ : Span4Mux_v
    port map (
            O => \N__2531\,
            I => \N__2528\
        );

    \I__233\ : Odrv4
    port map (
            O => \N__2528\,
            I => \A_c_18\
        );

    \I__232\ : InMux
    port map (
            O => \N__2525\,
            I => \N__2519\
        );

    \I__231\ : InMux
    port map (
            O => \N__2524\,
            I => \N__2519\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2519\,
            I => \N__2516\
        );

    \I__229\ : Sp12to4
    port map (
            O => \N__2516\,
            I => \N__2513\
        );

    \I__228\ : Span12Mux_v
    port map (
            O => \N__2513\,
            I => \N__2510\
        );

    \I__227\ : Odrv12
    port map (
            O => \N__2510\,
            I => \A_c_17\
        );

    \I__226\ : CascadeMux
    port map (
            O => \N__2507\,
            I => \U409_CIA.g0Z0Z_2_cascade_\
        );

    \I__225\ : ClkMux
    port map (
            O => \N__2504\,
            I => \N__2474\
        );

    \I__224\ : ClkMux
    port map (
            O => \N__2503\,
            I => \N__2474\
        );

    \I__223\ : ClkMux
    port map (
            O => \N__2502\,
            I => \N__2474\
        );

    \I__222\ : ClkMux
    port map (
            O => \N__2501\,
            I => \N__2474\
        );

    \I__221\ : ClkMux
    port map (
            O => \N__2500\,
            I => \N__2474\
        );

    \I__220\ : ClkMux
    port map (
            O => \N__2499\,
            I => \N__2474\
        );

    \I__219\ : ClkMux
    port map (
            O => \N__2498\,
            I => \N__2474\
        );

    \I__218\ : ClkMux
    port map (
            O => \N__2497\,
            I => \N__2474\
        );

    \I__217\ : ClkMux
    port map (
            O => \N__2496\,
            I => \N__2474\
        );

    \I__216\ : ClkMux
    port map (
            O => \N__2495\,
            I => \N__2474\
        );

    \I__215\ : GlobalMux
    port map (
            O => \N__2474\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.TACK_EN_iC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            I => \N__2504\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            I => \N__2503\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            I => \N__2502\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            I => \N__2498\
        );

    \INVU409_TRANSFER_ACK.CIA_ENABLED_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            I => \N__2495\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__2501\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__2500\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__2497\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            I => \N__2499\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            I => \N__2496\
        );

    \IN_MUX_bfv_11_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_5_0_\
        );

    \IN_MUX_bfv_11_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_11_6_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_13_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_7_0_\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2608\,
            in1 => \N__2889\,
            in2 => \N__2555\,
            in3 => \N__2524\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_11_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4384\,
            in1 => \N__4296\,
            in2 => \N__3020\,
            in3 => \N__2554\,
            lcout => \U409_CIA.g0Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_8_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__2525\,
            in1 => \N__2849\,
            in2 => \_gnd_net_\,
            in3 => \N__4468\,
            lcout => \U409_CIA.g0Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_2_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2684\,
            in2 => \_gnd_net_\,
            in3 => \N__2792\,
            lcout => OPEN,
            ltout => \U409_CIA.g0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_13_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2765\,
            in1 => \N__2816\,
            in2 => \N__2507\,
            in3 => \N__2738\,
            lcout => \U409_CIA.g0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_3_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__2764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2784\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__2842\,
            in1 => \N__2809\,
            in2 => \N__2852\,
            in3 => \N__2627\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2841\,
            in1 => \N__2808\,
            in2 => \N__2788\,
            in3 => \N__2763\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_10_LC_1_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__2708\,
            in1 => \N__6152\,
            in2 => \N__2654\,
            in3 => \N__2729\,
            lcout => \U409_CIA.g0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_1_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2706\,
            in1 => \N__2727\,
            in2 => \N__2653\,
            in3 => \N__2676\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_4_LC_1_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2728\,
            in1 => \N__2707\,
            in2 => \N__2683\,
            in3 => \N__2649\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.g0_14_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2890\,
            in1 => \N__2621\,
            in2 => \N__2615\,
            in3 => \N__2585\,
            lcout => \U409_CIA.g0Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_LC_3_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__2579\,
            in1 => \N__2933\,
            in2 => \_gnd_net_\,
            in3 => \N__2567\,
            lcout => \AUTOVECTORm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_0_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4282\,
            in2 => \_gnd_net_\,
            in3 => \N__3013\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACEm_3\,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEm_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_0_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4459\,
            in1 => \N__4366\,
            in2 => \N__2558\,
            in3 => \N__3037\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_1_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4365\,
            in1 => \N__2999\,
            in2 => \N__4292\,
            in3 => \N__3043\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_3_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4458\,
            in1 => \N__4281\,
            in2 => \N__3047\,
            in3 => \N__3000\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2978\,
            in1 => \N__2969\,
            in2 => \N__6151\,
            in3 => \N__2951\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__2924\,
            in1 => \N__4457\,
            in2 => \N__5658\,
            in3 => \N__6147\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACEm_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PORTSIZE_0_i_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__5644\,
            in1 => \N__4367\,
            in2 => \N__2912\,
            in3 => \N__3636\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.HIROM_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2897\,
            in1 => \N__4371\,
            in2 => \N__4460\,
            in3 => \N__2891\,
            lcout => \U409_ADDRESS_DECODE.HIROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3312\,
            in2 => \N__3299\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3154\,
            in2 => \_gnd_net_\,
            in3 => \N__2855\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3085\,
            in2 => \_gnd_net_\,
            in3 => \N__3074\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3118\,
            in2 => \_gnd_net_\,
            in3 => \N__3071\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3097\,
            in2 => \_gnd_net_\,
            in3 => \N__3068\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3250\,
            in2 => \_gnd_net_\,
            in3 => \N__3065\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3130\,
            in2 => \_gnd_net_\,
            in3 => \N__3062\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3142\,
            in2 => \_gnd_net_\,
            in3 => \N__3059\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__5127\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3211\,
            in2 => \_gnd_net_\,
            in3 => \N__3056\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3340\,
            in2 => \_gnd_net_\,
            in3 => \N__3053\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3407\,
            in2 => \_gnd_net_\,
            in3 => \N__3050\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3358\,
            in2 => \_gnd_net_\,
            in3 => \N__3182\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3193\,
            in2 => \_gnd_net_\,
            in3 => \N__3179\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3268\,
            in2 => \_gnd_net_\,
            in3 => \N__3176\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3229\,
            in2 => \_gnd_net_\,
            in3 => \N__3173\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3167\,
            in2 => \_gnd_net_\,
            in3 => \N__3170\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3166\,
            in1 => \N__3155\,
            in2 => \N__3319\,
            in3 => \N__3143\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3230\,
            in1 => \N__3131\,
            in2 => \N__3272\,
            in3 => \N__3119\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3501\,
            in1 => \N__3529\,
            in2 => \N__3107\,
            in3 => \N__3104\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__3098\,
            in1 => \N__3086\,
            in2 => \_gnd_net_\,
            in3 => \N__3296\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3365\,
            in1 => \N__3359\,
            in2 => \N__3347\,
            in3 => \N__3344\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3449\,
            in1 => \N__3500\,
            in2 => \N__3329\,
            in3 => \N__3326\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3297\,
            in1 => \_gnd_net_\,
            in2 => \N__3320\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__3448\,
            in1 => \N__3298\,
            in2 => \N__3544\,
            in3 => \N__3502\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5124\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3546\,
            in1 => \N__3497\,
            in2 => \N__3465\,
            in3 => \N__3278\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3406\,
            in1 => \N__3212\,
            in2 => \N__3257\,
            in3 => \N__3194\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3547\,
            in1 => \N__3460\,
            in2 => \N__3239\,
            in3 => \N__3236\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3548\,
            in1 => \N__3498\,
            in2 => \N__3466\,
            in3 => \N__3218\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3545\,
            in1 => \N__3496\,
            in2 => \N__3464\,
            in3 => \N__3200\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__3450\,
            in1 => \N__3559\,
            in2 => \N__3506\,
            in3 => \N__3543\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5122\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__3542\,
            in1 => \N__3499\,
            in2 => \N__3467\,
            in3 => \N__3416\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__3747\,
            in1 => \N__3392\,
            in2 => \N__3698\,
            in3 => \N__3780\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5947\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3391\,
            in1 => \N__3748\,
            in2 => \_gnd_net_\,
            in3 => \N__3693\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__5947\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__3863\,
            in1 => \N__3827\,
            in2 => \_gnd_net_\,
            in3 => \N__3688\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5948\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3373\,
            in2 => \N__3697\,
            in3 => \N__3802\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5948\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__3801\,
            in1 => \N__3847\,
            in2 => \N__3377\,
            in3 => \N__3692\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3C_net\,
            ce => 'H',
            sr => \N__5948\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIISJM1_2_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3919\,
            in1 => \N__3943\,
            in2 => \N__3983\,
            in3 => \N__3826\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3781\,
            in2 => \N__3380\,
            in3 => \N__3749\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5675\,
            in1 => \N__3637\,
            in2 => \_gnd_net_\,
            in3 => \N__4385\,
            lcout => \U409_ADDRESS_DECODE.un1_nREGSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nREGSPACE_i_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__3644\,
            in1 => \N__5674\,
            in2 => \_gnd_net_\,
            in3 => \N__4392\,
            lcout => \U409_ADDRESS_DECODE_un1_nREGSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4542\,
            in2 => \N__4739\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_5_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4558\,
            in2 => \_gnd_net_\,
            in3 => \N__3590\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4693\,
            in2 => \_gnd_net_\,
            in3 => \N__3587\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4750\,
            in2 => \_gnd_net_\,
            in3 => \N__3584\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4762\,
            in2 => \_gnd_net_\,
            in3 => \N__3581\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4504\,
            in2 => \_gnd_net_\,
            in3 => \N__3578\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4810\,
            in2 => \_gnd_net_\,
            in3 => \N__3575\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__5120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5146\,
            in2 => \_gnd_net_\,
            in3 => \N__3671\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4774\,
            in2 => \_gnd_net_\,
            in3 => \N__3668\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_11_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4828\,
            in2 => \_gnd_net_\,
            in3 => \N__3665\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4708\,
            in2 => \_gnd_net_\,
            in3 => \N__3662\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4570\,
            in2 => \_gnd_net_\,
            in3 => \N__3659\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4840\,
            in2 => \_gnd_net_\,
            in3 => \N__3656\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4672\,
            in2 => \_gnd_net_\,
            in3 => \N__3653\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4799\,
            in3 => \N__3650\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4529\,
            in2 => \_gnd_net_\,
            in3 => \N__3647\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LOWROM_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4301\,
            in1 => \N__4394\,
            in2 => \N__5600\,
            in3 => \N__4472\,
            lcout => \U409_ADDRESS_DECODE.LOWROMZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5273\,
            in1 => \N__5195\,
            in2 => \N__3872\,
            in3 => \N__5236\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5126\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_3_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3982\,
            in1 => \N__3920\,
            in2 => \_gnd_net_\,
            in3 => \N__3944\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIV9KM1_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__3746\,
            in1 => \N__3824\,
            in2 => \N__3782\,
            in3 => \N__3843\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_6_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3797\,
            in1 => \N__3969\,
            in2 => \N__3713\,
            in3 => \N__3854\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3940\,
            in2 => \_gnd_net_\,
            in3 => \N__3917\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIS6KM1_7_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__3848\,
            in1 => \N__3825\,
            in2 => \N__3803\,
            in3 => \N__3968\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_5_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3776\,
            in1 => \N__3745\,
            in2 => \N__3716\,
            in3 => \N__3709\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIRGA77_5_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__4151\,
            in1 => \N__4110\,
            in2 => \N__3701\,
            in3 => \N__3891\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__3971\,
            in1 => \_gnd_net_\,
            in2 => \N__3986\,
            in3 => \N__3941\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5943\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110011"
        )
    port map (
            in0 => \N__4150\,
            in1 => \N__3970\,
            in2 => \N__4114\,
            in3 => \N__3892\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5943\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__3972\,
            in1 => \N__3918\,
            in2 => \_gnd_net_\,
            in3 => \N__3942\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__5943\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__4867\,
            in1 => \N__3899\,
            in2 => \_gnd_net_\,
            in3 => \N__3893\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__5936\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_am_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000111"
        )
    port map (
            in0 => \N__4903\,
            in1 => \N__4923\,
            in2 => \N__4976\,
            in3 => \N__4480\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.m9_am_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__6106\,
            in1 => \N__4954\,
            in2 => \N__3878\,
            in3 => \N__4487\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m11_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001010111"
        )
    port map (
            in0 => \N__4952\,
            in1 => \N__4924\,
            in2 => \N__4907\,
            in3 => \N__4481\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.i6_mux_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__6107\,
            in1 => \N__4974\,
            in2 => \N__3875\,
            in3 => \N__4953\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIIJ4U_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4951\,
            in1 => \N__4877\,
            in2 => \N__4105\,
            in3 => \N__4891\,
            lcout => \U409_TRANSFER_ACK.N_105\,
            ltout => \U409_TRANSFER_ACK.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m9_bm_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101000111"
        )
    port map (
            in0 => \N__4922\,
            in1 => \N__4973\,
            in2 => \N__4490\,
            in3 => \N__4902\,
            lcout => \U409_TRANSFER_ACK.m9_bm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_ns_1_0__m3_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4876\,
            in2 => \_gnd_net_\,
            in3 => \N__4890\,
            lcout => \U409_TRANSFER_ACK.N_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un5_nRAMSPACE_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4464\,
            in1 => \N__4393\,
            in2 => \_gnd_net_\,
            in3 => \N__4300\,
            lcout => \U409_ADDRESS_DECODE.un5_nRAMSPACEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__5683\,
            in1 => \N__4228\,
            in2 => \N__4214\,
            in3 => \N__6108\,
            lcout => \ROMENm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMENm_i_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__6109\,
            in1 => \N__5676\,
            in2 => \N__4232\,
            in3 => \N__4213\,
            lcout => \ROMENm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER15_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__4166\,
            in1 => \N__4138\,
            in2 => \N__4106\,
            in3 => \N__4049\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS0_i_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__4025\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4660\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nCIACS1_i_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4646\,
            in2 => \_gnd_net_\,
            in3 => \N__4661\,
            lcout => \U409_ADDRESS_DECODE_un1_nCIACS1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_nRAMSPACE_i_LC_12_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__5711\,
            in1 => \N__5673\,
            in2 => \_gnd_net_\,
            in3 => \N__5589\,
            lcout => \U409_ADDRESS_DECODE_un1_nRAMSPACE_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__4546\,
            in1 => \N__4738\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5233\,
            in1 => \N__5266\,
            in2 => \N__5202\,
            in3 => \N__4601\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__5265\,
            in1 => \N__5235\,
            in2 => \N__5204\,
            in3 => \N__4582\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4571\,
            in1 => \N__4559\,
            in2 => \N__4547\,
            in3 => \N__4528\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__5264\,
            in1 => \N__5234\,
            in2 => \N__4517\,
            in3 => \N__5192\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5147\,
            in1 => \N__4775\,
            in2 => \N__4508\,
            in3 => \N__4673\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__4737\,
            in1 => \N__5232\,
            in2 => \N__4493\,
            in3 => \N__5269\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4841\,
            in1 => \N__4829\,
            in2 => \N__4817\,
            in3 => \N__4798\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5193\,
            in1 => \N__5268\,
            in2 => \N__4784\,
            in3 => \N__4781\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4763\,
            in1 => \N__4751\,
            in2 => \_gnd_net_\,
            in3 => \N__4736\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4715\,
            in1 => \N__4709\,
            in2 => \N__4697\,
            in3 => \N__4694\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5231\,
            in1 => \N__5194\,
            in2 => \N__4682\,
            in3 => \N__4679\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_RNIFVN95_0_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__4990\,
            in1 => \N__5071\,
            in2 => \N__5054\,
            in3 => \N__5029\,
            lcout => \CIA_ENABLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_HOLD_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__5070\,
            in1 => \N__5049\,
            in2 => \N__5030\,
            in3 => \N__4989\,
            lcout => \U409_CIA.CIA_HOLDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000100010"
        )
    port map (
            in0 => \N__5866\,
            in1 => \N__5482\,
            in2 => \_gnd_net_\,
            in3 => \N__5444\,
            lcout => OPEN,
            ltout => \U409_CIA.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101010101010"
        )
    port map (
            in0 => \N__5048\,
            in1 => \N__5867\,
            in2 => \N__4649\,
            in3 => \N__5762\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5385\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__5078\,
            in1 => \N__5053\,
            in2 => \N__5025\,
            in3 => \N__4994\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_ENABLED_0C_net\,
            ce => 'H',
            sr => \N__5742\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5410\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100011101000000"
        )
    port map (
            in0 => \N__4975\,
            in1 => \N__4955\,
            in2 => \N__4934\,
            in3 => \N__4853\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4925\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4892\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_0C_net\,
            ce => 'H',
            sr => \N__5749\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIHST5_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4868\,
            in2 => \_gnd_net_\,
            in3 => \N__4852\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110100000"
        )
    port map (
            in0 => \N__5348\,
            in1 => \_gnd_net_\,
            in2 => \N__5306\,
            in3 => \N__5327\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111110"
        )
    port map (
            in0 => \N__5325\,
            in1 => \N__5304\,
            in2 => \N__5368\,
            in3 => \N__5346\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100101010"
        )
    port map (
            in0 => \N__5279\,
            in1 => \N__5354\,
            in2 => \N__5369\,
            in3 => \N__5528\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111001100"
        )
    port map (
            in0 => \N__5326\,
            in1 => \N__5300\,
            in2 => \_gnd_net_\,
            in3 => \N__5347\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__5750\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5323\,
            in1 => \N__5344\,
            in2 => \_gnd_net_\,
            in3 => \N__5296\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__5345\,
            in1 => \N__5324\,
            in2 => \N__5305\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__5267\,
            in1 => \N__5237\,
            in2 => \N__5203\,
            in3 => \N__5156\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5118\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5439\,
            in2 => \N__5483\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_13_7_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5780\,
            in2 => \_gnd_net_\,
            in3 => \N__5087\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__5386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5861\,
            in2 => \_gnd_net_\,
            in3 => \N__5084\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5803\,
            in2 => \_gnd_net_\,
            in3 => \N__5081\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__5386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNO_0_5_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5829\,
            in2 => \_gnd_net_\,
            in3 => \N__5507\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT_RNO_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__5862\,
            in1 => \N__5501\,
            in2 => \N__5504\,
            in3 => \N__5477\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__5440\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5478\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5386\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIKSMD1_5_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5442\,
            in1 => \N__5782\,
            in2 => \N__5831\,
            in3 => \N__5804\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010011001100110"
        )
    port map (
            in0 => \N__5865\,
            in1 => \N__5495\,
            in2 => \N__5489\,
            in3 => \N__5481\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_2_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5863\,
            in1 => \N__5479\,
            in2 => \_gnd_net_\,
            in3 => \N__5441\,
            lcout => OPEN,
            ltout => \U409_CIA.N_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_0_LC_13_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5403\,
            in2 => \N__5486\,
            in3 => \N__5761\,
            lcout => OPEN,
            ltout => \U409_CIA.CLKCIAZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__5837\,
            in1 => \N__5480\,
            in2 => \N__5447\,
            in3 => \N__5443\,
            lcout => \CLKCIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5384\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLKCIA_RNO_1_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5802\,
            in1 => \N__5783\,
            in2 => \N__5830\,
            in3 => \N__5864\,
            lcout => \U409_CIA.CLKCIA6_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIH7921_5_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__5822\,
            in1 => \N__5801\,
            in2 => \_gnd_net_\,
            in3 => \N__5781\,
            lcout => \U409_CIA.CLKCIA8_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6089\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AGNUS_SPACE_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010101"
        )
    port map (
            in0 => \N__5723\,
            in1 => \N__5710\,
            in2 => \N__5687\,
            in3 => \N__5593\,
            lcout => \nBUFEN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__6185\,
            in1 => \_gnd_net_\,
            in2 => \N__6125\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011101010"
        )
    port map (
            in0 => \N__5539\,
            in1 => \N__6199\,
            in2 => \N__6126\,
            in3 => \N__6173\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNIURL11_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__6183\,
            in1 => \N__5527\,
            in2 => \N__6200\,
            in3 => \N__5516\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER_ns_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5510\,
            in3 => \N__6112\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_RNO_0_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__6116\,
            in1 => \N__6198\,
            in2 => \_gnd_net_\,
            in3 => \N__6184\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER_nss_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_i_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__6110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6172\,
            lcout => \TACK_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_EN_iC_net\,
            ce => \N__6161\,
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__6111\,
            in1 => \N__5983\,
            in2 => \_gnd_net_\,
            in3 => \N__5969\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \TACKn_iobuf_RNO_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_365_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 13 2025 12:13:37

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U400_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U400_TOP
entity U400_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    MA : out std_logic_vector(12 downto 0);
    A : in std_logic_vector(31 downto 0);
    LBENn : out std_logic;
    CS0n : out std_logic;
    UUBEn : out std_logic;
    TAn : out std_logic;
    CLK40 : in std_logic;
    RnW : in std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    WEn : out std_logic;
    LLBEn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    RASn : out std_logic;
    CS1n : out std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic);
end U400_TOP;

-- Architecture of U400_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U400_TOP is

signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7440\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7431\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7377\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7368\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7350\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7341\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7332\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7323\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7161\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7134\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7098\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7071\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7035\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6663\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6357\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6288\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5577\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5565\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5553\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5535\ : std_logic;
signal \N__5532\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5454\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5400\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5321\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5145\ : std_logic;
signal \N__5142\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5123\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5084\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5007\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5001\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4845\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4608\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4566\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4491\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4488\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4332\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4329\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4323\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4170\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4074\ : std_logic;
signal \N__4071\ : std_logic;
signal \N__4068\ : std_logic;
signal \N__4065\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3954\ : std_logic;
signal \N__3951\ : std_logic;
signal \N__3948\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3942\ : std_logic;
signal \N__3939\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3864\ : std_logic;
signal \N__3861\ : std_logic;
signal \N__3858\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3852\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3825\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3801\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3790\ : std_logic;
signal \N__3787\ : std_logic;
signal \N__3784\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3772\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3706\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3684\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3657\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3634\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3591\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3567\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3497\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3480\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3471\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3465\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3435\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3303\ : std_logic;
signal \N__3300\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3270\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3225\ : std_logic;
signal \N__3222\ : std_logic;
signal \N__3219\ : std_logic;
signal \N__3216\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3186\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3166\ : std_logic;
signal \N__3163\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3115\ : std_logic;
signal \N__3112\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3094\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3087\ : std_logic;
signal \N__3084\ : std_logic;
signal \N__3081\ : std_logic;
signal \N__3078\ : std_logic;
signal \N__3075\ : std_logic;
signal \N__3072\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3039\ : std_logic;
signal \N__3036\ : std_logic;
signal \N__3033\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3006\ : std_logic;
signal \N__3003\ : std_logic;
signal \N__3000\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2977\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2971\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2940\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2937\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2910\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2904\ : std_logic;
signal \N__2901\ : std_logic;
signal \N__2898\ : std_logic;
signal \N__2895\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2881\ : std_logic;
signal \N__2878\ : std_logic;
signal \N__2869\ : std_logic;
signal \N__2868\ : std_logic;
signal \N__2865\ : std_logic;
signal \N__2862\ : std_logic;
signal \N__2857\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2848\ : std_logic;
signal \N__2845\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2812\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2803\ : std_logic;
signal \N__2800\ : std_logic;
signal \N__2797\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2743\ : std_logic;
signal \N__2740\ : std_logic;
signal \N__2737\ : std_logic;
signal \N__2734\ : std_logic;
signal \N__2731\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2722\ : std_logic;
signal \N__2719\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2707\ : std_logic;
signal \CLK40_ibuf_gb_io_gb_input\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\ : std_logic;
signal \U400_SDRAM.CO1\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_31\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_27\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER23_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa\ : std_logic;
signal \U400_SDRAM.TA_COUNTER23\ : std_logic;
signal \U400_SDRAM.TA_COUNTER27\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\ : std_logic;
signal \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\ : std_logic;
signal \U400_SDRAM.BURSTZ0\ : std_logic;
signal \INVU400_SDRAM.BURSTC_net\ : std_logic;
signal \U400_SDRAM.TACKZ0\ : std_logic;
signal \INVU400_SDRAM.TACKC_net\ : std_logic;
signal \A_c_22\ : std_logic;
signal \BANK1_c\ : std_logic;
signal \A_c_21\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \INVU400_SDRAM.BANK1C_net\ : std_logic;
signal \RASn_c\ : std_logic;
signal \INVU400_SDRAM.RASnC_net\ : std_logic;
signal \U400_SDRAM.N_299_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_2C_net\ : std_logic;
signal \U400_SDRAM.N_52\ : std_logic;
signal \U400_SDRAM.N_295_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_300_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_0C_net\ : std_logic;
signal \U400_SDRAM.N_110_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_55_cascade_\ : std_logic;
signal \U400_SDRAM.N_105_cascade_\ : std_logic;
signal \U400_SDRAM.N_68\ : std_logic;
signal \U400_SDRAM.N_62_cascade_\ : std_logic;
signal \U400_SDRAM.N_39_cascade_\ : std_logic;
signal \U400_SDRAM.N_62\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U400_SDRAM.N_41_cascade_\ : std_logic;
signal \INVU400_SDRAM.CS0_ENC_net\ : std_logic;
signal \U400_SDRAM.N_57_cascade_\ : std_logic;
signal \U400_SDRAM.N_46\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_266_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD12\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD12_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_0\ : std_logic;
signal \U400_SDRAM.CS0_ENZ0\ : std_logic;
signal \CS0n_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \CASn_c\ : std_logic;
signal \INVU400_SDRAM.CS0nC_net\ : std_logic;
signal \U400_SDRAM.CS1_ENZ0\ : std_logic;
signal \CS1n_c\ : std_logic;
signal \INVU400_SDRAM.CS1nC_net\ : std_logic;
signal \A_c_9\ : std_logic;
signal \A_c_17\ : std_logic;
signal \MA_c_7\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_7C_net\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_16\ : std_logic;
signal \MA_c_6\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_6C_net\ : std_logic;
signal \bfn_5_4_0_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1\ : std_logic;
signal \U400_SDRAM.N_111\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U400_SDRAM.un3_RAM_CYCLE_START_cascade_\ : std_logic;
signal \U400_SDRAM.RAM_CYCLE_STARTZ0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.N_54_cascade_\ : std_logic;
signal \U400_SDRAM.N_57\ : std_logic;
signal \U400_SDRAM.N_51\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_0\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\ : std_logic;
signal \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\ : std_logic;
signal \INVU400_SDRAM.REFRESH_COUNTER_2C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\ : std_logic;
signal \A_c_24\ : std_logic;
signal \A_c_18\ : std_logic;
signal \MA_c_8\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_8C_net\ : std_logic;
signal \A_c_19\ : std_logic;
signal \MA_c_9\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_9C_net\ : std_logic;
signal \U400_SDRAM.N_110\ : std_logic;
signal \RnW_c\ : std_logic;
signal \INVU400_SDRAM.WRITE_CYCLEC_net\ : std_logic;
signal \U400_SDRAM.TA_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.TA_EN11_m\ : std_logic;
signal \U400_SDRAM.un1_TA_COUNTER26_2_0\ : std_logic;
signal \TA_OUT\ : std_logic;
signal \CLK40_c_g\ : std_logic;
signal \U400_SDRAM.N_105\ : std_logic;
signal \U400_SDRAM.N_59\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_\ : std_logic;
signal \U400_SDRAM.N_84\ : std_logic;
signal \U400_SDRAM.RAM_CYCLEZ0\ : std_logic;
signal \INVU400_SDRAM.RAM_CYCLEC_net\ : std_logic;
signal \U400_SDRAM.N_30_2_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0\ : std_logic;
signal \U400_SDRAM.N_30_2\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER44_5_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_117\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER42\ : std_logic;
signal \U400_SDRAM.un1_SDRAM_COUNTER44_0\ : std_logic;
signal \U400_SDRAM.TACK_4_m\ : std_logic;
signal \U400_SDRAM.TACK_7_0\ : std_logic;
signal \U400_SDRAM.N_56\ : std_logic;
signal \U400_SDRAM.N_56_cascade_\ : std_logic;
signal \U400_SDRAM.N_108\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_94_1\ : std_logic;
signal \U400_SDRAM.N_275_cascade_\ : std_logic;
signal \U400_SDRAM.N_54\ : std_logic;
signal \U400_SDRAM.N_276\ : std_logic;
signal \A_c_26\ : std_logic;
signal \MA_c_12\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_12C_net\ : std_logic;
signal \A_c_20\ : std_logic;
signal \MA_c_10\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_10C_net\ : std_logic;
signal \U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_\ : std_logic;
signal \U400_BYTE_ENABLE_un1_LLBEn_i\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0\ : std_logic;
signal \U400_SDRAM.N_321_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_322_0\ : std_logic;
signal \U400_SDRAM.WRITE_CYCLEZ0\ : std_logic;
signal \U400_SDRAM.N_320_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U400_SDRAM.N_88\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_3\ : std_logic;
signal \U400_SDRAM.N_303_0_i\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_5_sqmuxa\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \INVU400_SDRAM.SDRAM_COUNTER_0C_net\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\ : std_logic;
signal \U400_SDRAM.N_66\ : std_logic;
signal \U400_SDRAM.N_55\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0\ : std_logic;
signal \U400_SDRAM.REFRESH_COUNTERZ0Z_8\ : std_logic;
signal \U400_SDRAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U400_SDRAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0\ : std_logic;
signal \U400_SDRAM.N_299_2\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_\ : std_logic;
signal \U400_SDRAM.N_266_0\ : std_logic;
signal \U400_SDRAM.N_270\ : std_logic;
signal \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_\ : std_logic;
signal \U400_SDRAM.N_43\ : std_logic;
signal \INVU400_SDRAM.SDRAM_CMD_1C_net\ : std_logic;
signal \A_c_25\ : std_logic;
signal \MA_c_11\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_11C_net\ : std_logic;
signal \U400_BYTE_ENABLE_un1_UMBEn_i\ : std_logic;
signal \U400_BYTE_ENABLE_un1_LMBEn_i\ : std_logic;
signal \RAM_SPACEm\ : std_logic;
signal \U400_BYTE_ENABLE_un1_UUBEn_i\ : std_logic;
signal \A_c_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U400_BYTE_ENABLE.un2_UMBEn_0_0\ : std_logic;
signal \U400_BYTE_ENABLE.LW_TRANS_0\ : std_logic;
signal \U400_ADDRESS_DECODE_RAM_SPACE_3\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_28\ : std_logic;
signal \RAM_SPACEm_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \U400_SDRAM.BURSTZ0Z8\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_5\ : std_logic;
signal \MA_c_5\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_5C_net\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_13\ : std_logic;
signal \MA_c_3\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_3C_net\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_14\ : std_logic;
signal \MA_c_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_10\ : std_logic;
signal \MA_c_0\ : std_logic;
signal \A_c_11\ : std_logic;
signal \U400_SDRAM.MA_5_iv_0_1\ : std_logic;
signal \MA_c_1\ : std_logic;
signal \U400_SDRAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U400_SDRAM.MA19\ : std_logic;
signal \MA_c_2\ : std_logic;
signal \INVU400_SDRAM.MA_nesr_4C_net\ : std_logic;
signal \U400_SDRAM.un1_MA20_0_i_0\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \TA_EN_i_ess\ : std_logic;
signal \N_474_i\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \MA_wire\ : std_logic_vector(12 downto 0);
signal \A_wire\ : std_logic_vector(31 downto 0);
signal \CASn_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \UUBEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \LLBEn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \TAn_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CS1n_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CS0n_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CLK40_wire\ : std_logic;

begin
    MA <= \MA_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    BANK1 <= \BANK1_wire\;
    UUBEn <= \UUBEn_wire\;
    \SIZ_wire\ <= SIZ;
    LLBEn <= \LLBEn_wire\;
    \TSn_wire\ <= TSn;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    \RESETn_wire\ <= RESETn;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    TAn <= \TAn_wire\;
    LBENn <= \LBENn_wire\;
    CS1n <= \CS1n_wire\;
    WEn <= \WEn_wire\;
    \RnW_wire\ <= RnW;
    CS0n <= \CS0n_wire\;
    LMBEn <= \LMBEn_wire\;
    \CLK40_wire\ <= CLK40;

    \MA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7451\,
            DIN => \N__7450\,
            DOUT => \N__7449\,
            PACKAGEPIN => \MA_wire\(7)
        );

    \MA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7451\,
            PADOUT => \N__7450\,
            PADIN => \N__7449\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3400\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7442\,
            DIN => \N__7441\,
            DOUT => \N__7440\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7442\,
            PADOUT => \N__7441\,
            PADIN => \N__7440\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7433\,
            DIN => \N__7432\,
            DOUT => \N__7431\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7433\,
            PADOUT => \N__7432\,
            PADIN => \N__7431\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3238\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7424\,
            DIN => \N__7423\,
            DOUT => \N__7422\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7424\,
            PADOUT => \N__7423\,
            PADIN => \N__7422\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7415\,
            DIN => \N__7414\,
            DOUT => \N__7413\,
            PACKAGEPIN => \MA_wire\(8)
        );

    \MA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7415\,
            PADOUT => \N__7414\,
            PADIN => \N__7413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3736\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7406\,
            DIN => \N__7405\,
            DOUT => \N__7404\,
            PACKAGEPIN => \MA_wire\(10)
        );

    \MA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7406\,
            PADOUT => \N__7405\,
            PADIN => \N__7404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7397\,
            DIN => \N__7396\,
            DOUT => \N__7395\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7397\,
            PADOUT => \N__7396\,
            PADIN => \N__7395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7388\,
            DIN => \N__7387\,
            DOUT => \N__7386\,
            PACKAGEPIN => \MA_wire\(2)
        );

    \MA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7388\,
            PADOUT => \N__7387\,
            PADIN => \N__7386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6607\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7379\,
            DIN => \N__7378\,
            DOUT => \N__7377\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7379\,
            PADOUT => \N__7378\,
            PADIN => \N__7377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7370\,
            DIN => \N__7369\,
            DOUT => \N__7368\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7370\,
            PADOUT => \N__7369\,
            PADIN => \N__7368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7361\,
            DIN => \N__7360\,
            DOUT => \N__7359\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7361\,
            PADOUT => \N__7360\,
            PADIN => \N__7359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5824\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7352\,
            DIN => \N__7351\,
            DOUT => \N__7350\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7352\,
            PADOUT => \N__7351\,
            PADIN => \N__7350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7343\,
            DIN => \N__7342\,
            DOUT => \N__7341\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7343\,
            PADOUT => \N__7342\,
            PADIN => \N__7341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7334\,
            DIN => \N__7333\,
            DOUT => \N__7332\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7334\,
            PADOUT => \N__7333\,
            PADIN => \N__7332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7325\,
            DIN => \N__7324\,
            DOUT => \N__7323\,
            PACKAGEPIN => \MA_wire\(12)
        );

    \MA_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7325\,
            PADOUT => \N__7324\,
            PADIN => \N__7323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4267\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7316\,
            DIN => \N__7315\,
            DOUT => \N__7314\,
            PACKAGEPIN => \MA_wire\(1)
        );

    \MA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7316\,
            PADOUT => \N__7315\,
            PADIN => \N__7314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7307\,
            DIN => \N__7306\,
            DOUT => \N__7305\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7307\,
            PADOUT => \N__7306\,
            PADIN => \N__7305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7298\,
            DIN => \N__7297\,
            DOUT => \N__7296\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7298\,
            PADOUT => \N__7297\,
            PADIN => \N__7296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7289\,
            DIN => \N__7288\,
            DOUT => \N__7287\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7289\,
            PADOUT => \N__7288\,
            PADIN => \N__7287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7280\,
            DIN => \N__7279\,
            DOUT => \N__7278\,
            PACKAGEPIN => \MA_wire\(4)
        );

    \MA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7280\,
            PADOUT => \N__7279\,
            PADIN => \N__7278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5992\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7271\,
            DIN => \N__7270\,
            DOUT => \N__7269\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7271\,
            PADOUT => \N__7270\,
            PADIN => \N__7269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7262\,
            DIN => \N__7261\,
            DOUT => \N__7260\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7262\,
            PADOUT => \N__7261\,
            PADIN => \N__7260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7253\,
            DIN => \N__7252\,
            DOUT => \N__7251\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7253\,
            PADOUT => \N__7252\,
            PADIN => \N__7251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4522\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7244\,
            DIN => \N__7243\,
            DOUT => \N__7242\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7244\,
            PADOUT => \N__7243\,
            PADIN => \N__7242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7235\,
            DIN => \N__7234\,
            DOUT => \N__7233\,
            PACKAGEPIN => \MA_wire\(9)
        );

    \MA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7235\,
            PADOUT => \N__7234\,
            PADIN => \N__7233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3709\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7226\,
            DIN => \N__7225\,
            DOUT => \N__7224\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7226\,
            PADOUT => \N__7225\,
            PADIN => \N__7224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5863\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7217\,
            DIN => \N__7216\,
            DOUT => \N__7215\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7217\,
            PADOUT => \N__7216\,
            PADIN => \N__7215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7208\,
            DIN => \N__7207\,
            DOUT => \N__7206\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7208\,
            PADOUT => \N__7207\,
            PADIN => \N__7206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7199\,
            DIN => \N__7198\,
            DOUT => \N__7197\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7199\,
            PADOUT => \N__7198\,
            PADIN => \N__7197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2767\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7190\,
            DIN => \N__7189\,
            DOUT => \N__7188\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7190\,
            PADOUT => \N__7189\,
            PADIN => \N__7188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7181\,
            DIN => \N__7180\,
            DOUT => \N__7179\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7181\,
            PADOUT => \N__7180\,
            PADIN => \N__7179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7172\,
            DIN => \N__7171\,
            DOUT => \N__7170\,
            PACKAGEPIN => \MA_wire\(3)
        );

    \MA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7172\,
            PADOUT => \N__7171\,
            PADIN => \N__7170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7163\,
            DIN => \N__7162\,
            DOUT => \N__7161\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7163\,
            PADOUT => \N__7162\,
            PADIN => \N__7161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7154\,
            DIN => \N__7153\,
            DOUT => \N__7152\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7154\,
            PADOUT => \N__7153\,
            PADIN => \N__7152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7145\,
            DIN => \N__7144\,
            DOUT => \N__7143\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7145\,
            PADOUT => \N__7144\,
            PADIN => \N__7143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7136\,
            DIN => \N__7135\,
            DOUT => \N__7134\,
            PACKAGEPIN => \MA_wire\(6)
        );

    \MA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7136\,
            PADOUT => \N__7135\,
            PADIN => \N__7134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7127\,
            DIN => \N__7126\,
            DOUT => \N__7125\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7127\,
            PADOUT => \N__7126\,
            PADIN => \N__7125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7118\,
            DIN => \N__7117\,
            DOUT => \N__7116\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7118\,
            PADOUT => \N__7117\,
            PADIN => \N__7116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7109\,
            DIN => \N__7108\,
            DOUT => \N__7107\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7109\,
            PADOUT => \N__7108\,
            PADIN => \N__7107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7100\,
            DIN => \N__7099\,
            DOUT => \N__7098\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7100\,
            PADOUT => \N__7099\,
            PADIN => \N__7098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7091\,
            DIN => \N__7090\,
            DOUT => \N__7089\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7091\,
            PADOUT => \N__7090\,
            PADIN => \N__7089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7082\,
            DIN => \N__7081\,
            DOUT => \N__7080\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7082\,
            PADOUT => \N__7081\,
            PADIN => \N__7080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3013\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7073\,
            DIN => \N__7072\,
            DOUT => \N__7071\,
            PACKAGEPIN => \MA_wire\(11)
        );

    \MA_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7073\,
            PADOUT => \N__7072\,
            PADIN => \N__7071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5872\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7064\,
            DIN => \N__7063\,
            DOUT => \N__7062\,
            PACKAGEPIN => \TAn_wire\
        );

    \TAn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7064\,
            PADOUT => \N__7063\,
            PADIN => \N__7062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__6412\,
            DIN0 => OPEN,
            DOUT0 => \N__4084\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7055\,
            DIN => \N__7054\,
            DOUT => \N__7053\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7055\,
            PADOUT => \N__7054\,
            PADIN => \N__7053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7046\,
            DIN => \N__7045\,
            DOUT => \N__7044\,
            PACKAGEPIN => \MA_wire\(5)
        );

    \MA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7046\,
            PADOUT => \N__7045\,
            PADIN => \N__7044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6076\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7037\,
            DIN => \N__7036\,
            DOUT => \N__7035\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7037\,
            PADOUT => \N__7036\,
            PADIN => \N__7035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7028\,
            DIN => \N__7027\,
            DOUT => \N__7026\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7028\,
            PADOUT => \N__7027\,
            PADIN => \N__7026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LBENn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7019\,
            DIN => \N__7018\,
            DOUT => \N__7017\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7019\,
            PADOUT => \N__7018\,
            PADIN => \N__7017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5599\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7010\,
            DIN => \N__7009\,
            DOUT => \N__7008\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7010\,
            PADOUT => \N__7009\,
            PADIN => \N__7008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7001\,
            DIN => \N__7000\,
            DOUT => \N__6999\,
            PACKAGEPIN => \CS1n_wire\
        );

    \CS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7001\,
            PADOUT => \N__7000\,
            PADIN => \N__6999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3211\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6992\,
            DIN => \N__6991\,
            DOUT => \N__6990\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6992\,
            PADOUT => \N__6991\,
            PADIN => \N__6990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6983\,
            DIN => \N__6982\,
            DOUT => \N__6981\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6983\,
            PADOUT => \N__6982\,
            PADIN => \N__6981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6974\,
            DIN => \N__6973\,
            DOUT => \N__6972\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6974\,
            PADOUT => \N__6973\,
            PADIN => \N__6972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6965\,
            DIN => \N__6964\,
            DOUT => \N__6963\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6965\,
            PADOUT => \N__6964\,
            PADIN => \N__6963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6956\,
            DIN => \N__6955\,
            DOUT => \N__6954\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6956\,
            PADOUT => \N__6955\,
            PADIN => \N__6954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3247\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \MA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6947\,
            DIN => \N__6946\,
            DOUT => \N__6945\,
            PACKAGEPIN => \MA_wire\(0)
        );

    \MA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6947\,
            PADOUT => \N__6946\,
            PADIN => \N__6945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5950\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6938\,
            DIN => \N__6937\,
            DOUT => \N__6936\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6938\,
            PADOUT => \N__6937\,
            PADIN => \N__6936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6929\,
            DIN => \N__6928\,
            DOUT => \N__6927\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6929\,
            PADOUT => \N__6928\,
            PADIN => \N__6927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6920\,
            DIN => \N__6919\,
            DOUT => \N__6918\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6920\,
            PADOUT => \N__6919\,
            PADIN => \N__6918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6911\,
            DIN => \N__6910\,
            DOUT => \N__6909\,
            PACKAGEPIN => \CS0n_wire\
        );

    \CS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6911\,
            PADOUT => \N__6910\,
            PADIN => \N__6909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6902\,
            DIN => \N__6901\,
            DOUT => \N__6900\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6902\,
            PADOUT => \N__6901\,
            PADIN => \N__6900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6893\,
            DIN => \N__6892\,
            DOUT => \N__6891\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6893\,
            PADOUT => \N__6892\,
            PADIN => \N__6891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5854\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6884\,
            DIN => \N__6883\,
            DOUT => \N__6882\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6884\,
            PADOUT => \N__6883\,
            PADIN => \N__6882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6875\,
            DIN => \N__6874\,
            DOUT => \N__6873\,
            PACKAGEPIN => \CLK40_wire\
        );

    \CLK40_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6875\,
            PADOUT => \N__6874\,
            PADIN => \N__6873\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_ibuf_gb_io_gb_input\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1634\ : IoInMux
    port map (
            O => \N__6856\,
            I => \N__6853\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__6853\,
            I => \N__6850\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__6850\,
            I => \MA_c_1\
        );

    \I__1631\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6836\
        );

    \I__1630\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6827\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6827\
        );

    \I__1628\ : InMux
    port map (
            O => \N__6844\,
            I => \N__6827\
        );

    \I__1627\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6824\
        );

    \I__1626\ : InMux
    port map (
            O => \N__6842\,
            I => \N__6818\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6813\
        );

    \I__1624\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6813\
        );

    \I__1623\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6810\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__6836\,
            I => \N__6807\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6804\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6801\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__6827\,
            I => \N__6796\
        );

    \I__1618\ : LocalMux
    port map (
            O => \N__6824\,
            I => \N__6796\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6823\,
            I => \N__6793\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6790\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6787\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__6818\,
            I => \N__6780\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__6813\,
            I => \N__6780\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__6810\,
            I => \N__6780\
        );

    \I__1611\ : Span4Mux_v
    port map (
            O => \N__6807\,
            I => \N__6777\
        );

    \I__1610\ : LocalMux
    port map (
            O => \N__6804\,
            I => \N__6773\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__6801\,
            I => \N__6767\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__6796\,
            I => \N__6764\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__6793\,
            I => \N__6757\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__6790\,
            I => \N__6757\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__6787\,
            I => \N__6757\
        );

    \I__1604\ : Span4Mux_v
    port map (
            O => \N__6780\,
            I => \N__6754\
        );

    \I__1603\ : Sp12to4
    port map (
            O => \N__6777\,
            I => \N__6750\
        );

    \I__1602\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6747\
        );

    \I__1601\ : Span4Mux_s3_h
    port map (
            O => \N__6773\,
            I => \N__6744\
        );

    \I__1600\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6741\
        );

    \I__1599\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6738\
        );

    \I__1598\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6735\
        );

    \I__1597\ : Span4Mux_h
    port map (
            O => \N__6767\,
            I => \N__6732\
        );

    \I__1596\ : Span4Mux_h
    port map (
            O => \N__6764\,
            I => \N__6727\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__6757\,
            I => \N__6727\
        );

    \I__1594\ : Span4Mux_h
    port map (
            O => \N__6754\,
            I => \N__6724\
        );

    \I__1593\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6721\
        );

    \I__1592\ : Span12Mux_s8_h
    port map (
            O => \N__6750\,
            I => \N__6706\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__6747\,
            I => \N__6706\
        );

    \I__1590\ : Sp12to4
    port map (
            O => \N__6744\,
            I => \N__6706\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6741\,
            I => \N__6706\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6706\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__6735\,
            I => \N__6706\
        );

    \I__1586\ : Sp12to4
    port map (
            O => \N__6732\,
            I => \N__6706\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__6727\,
            I => \N__6703\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__6724\,
            I => \N__6700\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__6721\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1582\ : Odrv12
    port map (
            O => \N__6706\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1581\ : Odrv4
    port map (
            O => \N__6703\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1580\ : Odrv4
    port map (
            O => \N__6700\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_2\
        );

    \I__1579\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6688\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__6685\,
            I => \N__6682\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__6682\,
            I => \A_c_4\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__6679\,
            I => \N__6676\
        );

    \I__1574\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__6673\,
            I => \N__6670\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__6670\,
            I => \A_c_12\
        );

    \I__1571\ : InMux
    port map (
            O => \N__6667\,
            I => \N__6660\
        );

    \I__1570\ : InMux
    port map (
            O => \N__6666\,
            I => \N__6649\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6665\,
            I => \N__6649\
        );

    \I__1568\ : InMux
    port map (
            O => \N__6664\,
            I => \N__6649\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6663\,
            I => \N__6649\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6645\
        );

    \I__1565\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6642\
        );

    \I__1564\ : InMux
    port map (
            O => \N__6658\,
            I => \N__6639\
        );

    \I__1563\ : LocalMux
    port map (
            O => \N__6649\,
            I => \N__6635\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6648\,
            I => \N__6632\
        );

    \I__1561\ : Span12Mux_s4_v
    port map (
            O => \N__6645\,
            I => \N__6625\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6642\,
            I => \N__6625\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6639\,
            I => \N__6625\
        );

    \I__1558\ : InMux
    port map (
            O => \N__6638\,
            I => \N__6622\
        );

    \I__1557\ : Span4Mux_s2_v
    port map (
            O => \N__6635\,
            I => \N__6619\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__6632\,
            I => \N__6616\
        );

    \I__1555\ : Odrv12
    port map (
            O => \N__6625\,
            I => \U400_SDRAM.MA19\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6622\,
            I => \U400_SDRAM.MA19\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__6619\,
            I => \U400_SDRAM.MA19\
        );

    \I__1552\ : Odrv12
    port map (
            O => \N__6616\,
            I => \U400_SDRAM.MA19\
        );

    \I__1551\ : IoInMux
    port map (
            O => \N__6607\,
            I => \N__6604\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6601\
        );

    \I__1549\ : Odrv4
    port map (
            O => \N__6601\,
            I => \MA_c_2\
        );

    \I__1548\ : CEMux
    port map (
            O => \N__6598\,
            I => \N__6594\
        );

    \I__1547\ : CEMux
    port map (
            O => \N__6597\,
            I => \N__6589\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6594\,
            I => \N__6585\
        );

    \I__1545\ : CEMux
    port map (
            O => \N__6593\,
            I => \N__6582\
        );

    \I__1544\ : CEMux
    port map (
            O => \N__6592\,
            I => \N__6576\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6573\
        );

    \I__1542\ : CEMux
    port map (
            O => \N__6588\,
            I => \N__6570\
        );

    \I__1541\ : Span4Mux_s3_h
    port map (
            O => \N__6585\,
            I => \N__6564\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6582\,
            I => \N__6564\
        );

    \I__1539\ : CEMux
    port map (
            O => \N__6581\,
            I => \N__6561\
        );

    \I__1538\ : CEMux
    port map (
            O => \N__6580\,
            I => \N__6558\
        );

    \I__1537\ : CEMux
    port map (
            O => \N__6579\,
            I => \N__6555\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6576\,
            I => \N__6547\
        );

    \I__1535\ : Span4Mux_v
    port map (
            O => \N__6573\,
            I => \N__6547\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6570\,
            I => \N__6547\
        );

    \I__1533\ : CEMux
    port map (
            O => \N__6569\,
            I => \N__6544\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__6564\,
            I => \N__6535\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__6561\,
            I => \N__6535\
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6535\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6555\,
            I => \N__6535\
        );

    \I__1528\ : CEMux
    port map (
            O => \N__6554\,
            I => \N__6532\
        );

    \I__1527\ : Sp12to4
    port map (
            O => \N__6547\,
            I => \N__6527\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6544\,
            I => \N__6527\
        );

    \I__1525\ : Sp12to4
    port map (
            O => \N__6535\,
            I => \N__6522\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6532\,
            I => \N__6522\
        );

    \I__1523\ : Odrv12
    port map (
            O => \N__6527\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__6522\,
            I => \U400_SDRAM.un1_MA20_0_i_0\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6514\,
            I => \N__6510\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6513\,
            I => \N__6507\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6510\,
            I => \N__6497\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6483\
        );

    \I__1516\ : SRMux
    port map (
            O => \N__6506\,
            I => \N__6430\
        );

    \I__1515\ : SRMux
    port map (
            O => \N__6505\,
            I => \N__6430\
        );

    \I__1514\ : SRMux
    port map (
            O => \N__6504\,
            I => \N__6430\
        );

    \I__1513\ : SRMux
    port map (
            O => \N__6503\,
            I => \N__6430\
        );

    \I__1512\ : SRMux
    port map (
            O => \N__6502\,
            I => \N__6430\
        );

    \I__1511\ : SRMux
    port map (
            O => \N__6501\,
            I => \N__6430\
        );

    \I__1510\ : SRMux
    port map (
            O => \N__6500\,
            I => \N__6430\
        );

    \I__1509\ : Glb2LocalMux
    port map (
            O => \N__6497\,
            I => \N__6430\
        );

    \I__1508\ : SRMux
    port map (
            O => \N__6496\,
            I => \N__6430\
        );

    \I__1507\ : SRMux
    port map (
            O => \N__6495\,
            I => \N__6430\
        );

    \I__1506\ : SRMux
    port map (
            O => \N__6494\,
            I => \N__6430\
        );

    \I__1505\ : SRMux
    port map (
            O => \N__6493\,
            I => \N__6430\
        );

    \I__1504\ : SRMux
    port map (
            O => \N__6492\,
            I => \N__6430\
        );

    \I__1503\ : SRMux
    port map (
            O => \N__6491\,
            I => \N__6430\
        );

    \I__1502\ : SRMux
    port map (
            O => \N__6490\,
            I => \N__6430\
        );

    \I__1501\ : SRMux
    port map (
            O => \N__6489\,
            I => \N__6430\
        );

    \I__1500\ : SRMux
    port map (
            O => \N__6488\,
            I => \N__6430\
        );

    \I__1499\ : SRMux
    port map (
            O => \N__6487\,
            I => \N__6430\
        );

    \I__1498\ : SRMux
    port map (
            O => \N__6486\,
            I => \N__6430\
        );

    \I__1497\ : Glb2LocalMux
    port map (
            O => \N__6483\,
            I => \N__6430\
        );

    \I__1496\ : SRMux
    port map (
            O => \N__6482\,
            I => \N__6430\
        );

    \I__1495\ : SRMux
    port map (
            O => \N__6481\,
            I => \N__6430\
        );

    \I__1494\ : SRMux
    port map (
            O => \N__6480\,
            I => \N__6430\
        );

    \I__1493\ : SRMux
    port map (
            O => \N__6479\,
            I => \N__6430\
        );

    \I__1492\ : GlobalMux
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1491\ : gio2CtrlBuf
    port map (
            O => \N__6427\,
            I => \RESETn_c_i_g\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1488\ : Span12Mux_s6_h
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__1487\ : Odrv12
    port map (
            O => \N__6415\,
            I => \TA_EN_i_ess\
        );

    \I__1486\ : IoInMux
    port map (
            O => \N__6412\,
            I => \N__6409\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6409\,
            I => \N__6406\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__6406\,
            I => \N_474_i\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6397\
        );

    \I__1482\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6394\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6389\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6400\,
            I => \N__6389\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__6397\,
            I => \N__6385\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__6394\,
            I => \N__6382\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__6389\,
            I => \N__6379\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6376\
        );

    \I__1475\ : Sp12to4
    port map (
            O => \N__6385\,
            I => \N__6373\
        );

    \I__1474\ : Span4Mux_h
    port map (
            O => \N__6382\,
            I => \N__6370\
        );

    \I__1473\ : Span4Mux_h
    port map (
            O => \N__6379\,
            I => \N__6365\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6376\,
            I => \N__6365\
        );

    \I__1471\ : Span12Mux_s7_v
    port map (
            O => \N__6373\,
            I => \N__6362\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__6370\,
            I => \N__6357\
        );

    \I__1469\ : Span4Mux_v
    port map (
            O => \N__6365\,
            I => \N__6357\
        );

    \I__1468\ : Odrv12
    port map (
            O => \N__6362\,
            I => \SIZ_c_0\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__6357\,
            I => \SIZ_c_0\
        );

    \I__1466\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \N__6349\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6344\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__6348\,
            I => \N__6341\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__6347\,
            I => \N__6338\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6344\,
            I => \N__6335\
        );

    \I__1461\ : InMux
    port map (
            O => \N__6341\,
            I => \N__6332\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6329\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__6335\,
            I => \U400_SDRAM.BURSTZ0Z8\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6332\,
            I => \U400_SDRAM.BURSTZ0Z8\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6329\,
            I => \U400_SDRAM.BURSTZ0Z8\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1455\ : InMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1453\ : Odrv12
    port map (
            O => \N__6313\,
            I => \A_c_7\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \N__6302\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6309\,
            I => \N__6296\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6308\,
            I => \N__6296\
        );

    \I__1449\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6293\
        );

    \I__1448\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6289\
        );

    \I__1447\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6283\
        );

    \I__1446\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6280\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6277\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6274\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__6293\,
            I => \N__6271\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6292\,
            I => \N__6268\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6289\,
            I => \N__6265\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6288\,
            I => \N__6262\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6287\,
            I => \N__6259\
        );

    \I__1438\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6256\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6283\,
            I => \N__6244\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__6280\,
            I => \N__6244\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6244\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__6274\,
            I => \N__6244\
        );

    \I__1433\ : Span4Mux_h
    port map (
            O => \N__6271\,
            I => \N__6244\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6268\,
            I => \N__6241\
        );

    \I__1431\ : Span4Mux_h
    port map (
            O => \N__6265\,
            I => \N__6232\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6232\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6232\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6232\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6255\,
            I => \N__6229\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__6244\,
            I => \N__6226\
        );

    \I__1425\ : Span4Mux_h
    port map (
            O => \N__6241\,
            I => \N__6221\
        );

    \I__1424\ : Span4Mux_v
    port map (
            O => \N__6232\,
            I => \N__6221\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6229\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1422\ : Odrv4
    port map (
            O => \N__6226\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__6221\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_1\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__6214\,
            I => \N__6211\
        );

    \I__1419\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1417\ : Span4Mux_h
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1416\ : Odrv4
    port map (
            O => \N__6202\,
            I => \A_c_3\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6189\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6189\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6184\
        );

    \I__1412\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6181\
        );

    \I__1411\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6178\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6175\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6189\,
            I => \N__6172\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6167\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__6187\,
            I => \N__6164\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__6184\,
            I => \N__6160\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6157\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__6178\,
            I => \N__6154\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__6175\,
            I => \N__6149\
        );

    \I__1402\ : Span4Mux_s3_v
    port map (
            O => \N__6172\,
            I => \N__6149\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6146\
        );

    \I__1400\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6143\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6140\
        );

    \I__1398\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6135\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6135\
        );

    \I__1396\ : Span4Mux_v
    port map (
            O => \N__6160\,
            I => \N__6132\
        );

    \I__1395\ : Span4Mux_s3_v
    port map (
            O => \N__6157\,
            I => \N__6123\
        );

    \I__1394\ : Span4Mux_h
    port map (
            O => \N__6154\,
            I => \N__6123\
        );

    \I__1393\ : Span4Mux_h
    port map (
            O => \N__6149\,
            I => \N__6123\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6146\,
            I => \N__6123\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6143\,
            I => \N__6117\
        );

    \I__1390\ : Span4Mux_h
    port map (
            O => \N__6140\,
            I => \N__6117\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__6135\,
            I => \N__6110\
        );

    \I__1388\ : Span4Mux_h
    port map (
            O => \N__6132\,
            I => \N__6110\
        );

    \I__1387\ : Span4Mux_v
    port map (
            O => \N__6123\,
            I => \N__6110\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6122\,
            I => \N__6107\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__6117\,
            I => \N__6104\
        );

    \I__1384\ : Span4Mux_v
    port map (
            O => \N__6110\,
            I => \N__6101\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6107\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1382\ : Odrv4
    port map (
            O => \N__6104\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__6101\,
            I => \U400_SDRAM.SDRAM_CMDZ0Z_0\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6091\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6091\,
            I => \N__6088\
        );

    \I__1378\ : IoSpan4Mux
    port map (
            O => \N__6088\,
            I => \N__6085\
        );

    \I__1377\ : Odrv4
    port map (
            O => \N__6085\,
            I => \A_c_15\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6079\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6079\,
            I => \U400_SDRAM.MA_5_iv_0_5\
        );

    \I__1374\ : IoInMux
    port map (
            O => \N__6076\,
            I => \N__6073\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6073\,
            I => \N__6070\
        );

    \I__1372\ : IoSpan4Mux
    port map (
            O => \N__6070\,
            I => \N__6067\
        );

    \I__1371\ : IoSpan4Mux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__6064\,
            I => \MA_c_5\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6061\,
            I => \N__6058\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6055\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__6055\,
            I => \A_c_5\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6046\,
            I => \N__6043\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__6043\,
            I => \N__6040\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6040\,
            I => \A_c_13\
        );

    \I__1361\ : IoInMux
    port map (
            O => \N__6037\,
            I => \N__6034\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__6034\,
            I => \N__6031\
        );

    \I__1359\ : IoSpan4Mux
    port map (
            O => \N__6031\,
            I => \N__6028\
        );

    \I__1358\ : Span4Mux_s3_h
    port map (
            O => \N__6028\,
            I => \N__6025\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__6025\,
            I => \N__6022\
        );

    \I__1356\ : Odrv4
    port map (
            O => \N__6022\,
            I => \MA_c_3\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6016\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__6016\,
            I => \N__6013\
        );

    \I__1353\ : Span4Mux_s3_v
    port map (
            O => \N__6013\,
            I => \N__6010\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__6010\,
            I => \A_c_6\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__6007\,
            I => \N__6004\
        );

    \I__1350\ : InMux
    port map (
            O => \N__6004\,
            I => \N__6001\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6001\,
            I => \N__5998\
        );

    \I__1348\ : IoSpan4Mux
    port map (
            O => \N__5998\,
            I => \N__5995\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__5995\,
            I => \A_c_14\
        );

    \I__1346\ : IoInMux
    port map (
            O => \N__5992\,
            I => \N__5989\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__5989\,
            I => \N__5986\
        );

    \I__1344\ : IoSpan4Mux
    port map (
            O => \N__5986\,
            I => \N__5983\
        );

    \I__1343\ : Span4Mux_s1_v
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1342\ : Span4Mux_h
    port map (
            O => \N__5980\,
            I => \N__5977\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__5977\,
            I => \MA_c_4\
        );

    \I__1340\ : InMux
    port map (
            O => \N__5974\,
            I => \N__5971\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__5971\,
            I => \N__5968\
        );

    \I__1338\ : Span4Mux_h
    port map (
            O => \N__5968\,
            I => \N__5965\
        );

    \I__1337\ : Odrv4
    port map (
            O => \N__5965\,
            I => \A_c_2\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__5962\,
            I => \N__5959\
        );

    \I__1335\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5956\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__5956\,
            I => \N__5953\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__5953\,
            I => \A_c_10\
        );

    \I__1332\ : IoInMux
    port map (
            O => \N__5950\,
            I => \N__5947\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__5947\,
            I => \N__5944\
        );

    \I__1330\ : Span4Mux_s1_v
    port map (
            O => \N__5944\,
            I => \N__5941\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__5941\,
            I => \MA_c_0\
        );

    \I__1328\ : InMux
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__5935\,
            I => \N__5932\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__5932\,
            I => \A_c_11\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__5926\,
            I => \U400_SDRAM.MA_5_iv_0_1\
        );

    \I__1323\ : InMux
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5920\,
            I => \N__5917\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__5917\,
            I => \U400_SDRAM.N_270\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_\
        );

    \I__1319\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__1317\ : Span4Mux_h
    port map (
            O => \N__5905\,
            I => \N__5900\
        );

    \I__1316\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5897\
        );

    \I__1315\ : InMux
    port map (
            O => \N__5903\,
            I => \N__5894\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__5900\,
            I => \U400_SDRAM.N_43\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__5897\,
            I => \U400_SDRAM.N_43\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5894\,
            I => \U400_SDRAM.N_43\
        );

    \I__1311\ : CascadeMux
    port map (
            O => \N__5887\,
            I => \N__5884\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5881\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__5881\,
            I => \N__5878\
        );

    \I__1308\ : Span12Mux_v
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__5875\,
            I => \A_c_25\
        );

    \I__1306\ : IoInMux
    port map (
            O => \N__5872\,
            I => \N__5869\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__1304\ : Odrv12
    port map (
            O => \N__5866\,
            I => \MA_c_11\
        );

    \I__1303\ : IoInMux
    port map (
            O => \N__5863\,
            I => \N__5860\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__5860\,
            I => \N__5857\
        );

    \I__1301\ : Odrv4
    port map (
            O => \N__5857\,
            I => \U400_BYTE_ENABLE_un1_UMBEn_i\
        );

    \I__1300\ : IoInMux
    port map (
            O => \N__5854\,
            I => \N__5851\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5848\
        );

    \I__1298\ : Span4Mux_s2_v
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__1297\ : Odrv4
    port map (
            O => \N__5845\,
            I => \U400_BYTE_ENABLE_un1_LMBEn_i\
        );

    \I__1296\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5832\
        );

    \I__1295\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5832\
        );

    \I__1294\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5832\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5829\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5832\,
            I => \RAM_SPACEm\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5829\,
            I => \RAM_SPACEm\
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__1288\ : Span12Mux_s2_v
    port map (
            O => \N__5818\,
            I => \N__5815\
        );

    \I__1287\ : Odrv12
    port map (
            O => \N__5815\,
            I => \U400_BYTE_ENABLE_un1_UUBEn_i\
        );

    \I__1286\ : InMux
    port map (
            O => \N__5812\,
            I => \N__5808\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__5811\,
            I => \N__5805\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5800\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5805\,
            I => \N__5795\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5804\,
            I => \N__5795\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5792\
        );

    \I__1280\ : Span4Mux_v
    port map (
            O => \N__5800\,
            I => \N__5789\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5795\,
            I => \N__5784\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5792\,
            I => \N__5784\
        );

    \I__1277\ : Sp12to4
    port map (
            O => \N__5789\,
            I => \N__5781\
        );

    \I__1276\ : Span4Mux_h
    port map (
            O => \N__5784\,
            I => \N__5778\
        );

    \I__1275\ : Span12Mux_s6_h
    port map (
            O => \N__5781\,
            I => \N__5773\
        );

    \I__1274\ : Sp12to4
    port map (
            O => \N__5778\,
            I => \N__5773\
        );

    \I__1273\ : Span12Mux_v
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__1272\ : Odrv12
    port map (
            O => \N__5770\,
            I => \A_c_0\
        );

    \I__1271\ : CascadeMux
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5752\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5752\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5752\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5749\
        );

    \I__1266\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5744\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5744\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5737\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5749\,
            I => \N__5737\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5737\
        );

    \I__1261\ : Sp12to4
    port map (
            O => \N__5737\,
            I => \N__5734\
        );

    \I__1260\ : Span12Mux_v
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__1259\ : Odrv12
    port map (
            O => \N__5731\,
            I => \A_c_1\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__5725\,
            I => \U400_BYTE_ENABLE.un2_UMBEn_0_0\
        );

    \I__1256\ : CascadeMux
    port map (
            O => \N__5722\,
            I => \N__5718\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5713\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5713\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__5713\,
            I => \U400_BYTE_ENABLE.LW_TRANS_0\
        );

    \I__1252\ : CascadeMux
    port map (
            O => \N__5710\,
            I => \N__5706\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5702\
        );

    \I__1250\ : InMux
    port map (
            O => \N__5706\,
            I => \N__5699\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5705\,
            I => \N__5696\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5702\,
            I => \N__5693\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5699\,
            I => \N__5690\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5687\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__5693\,
            I => \N__5684\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__5690\,
            I => \N__5681\
        );

    \I__1243\ : Span12Mux_v
    port map (
            O => \N__5687\,
            I => \N__5676\
        );

    \I__1242\ : Sp12to4
    port map (
            O => \N__5684\,
            I => \N__5676\
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__5681\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_3\
        );

    \I__1240\ : Odrv12
    port map (
            O => \N__5676\,
            I => \U400_ADDRESS_DECODE_RAM_SPACE_3\
        );

    \I__1239\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5666\
        );

    \I__1238\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5663\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5660\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5666\,
            I => \N__5657\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5663\,
            I => \N__5654\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__5660\,
            I => \N__5651\
        );

    \I__1233\ : Span4Mux_h
    port map (
            O => \N__5657\,
            I => \N__5648\
        );

    \I__1232\ : Span4Mux_v
    port map (
            O => \N__5654\,
            I => \N__5643\
        );

    \I__1231\ : Span4Mux_h
    port map (
            O => \N__5651\,
            I => \N__5643\
        );

    \I__1230\ : Span4Mux_h
    port map (
            O => \N__5648\,
            I => \N__5640\
        );

    \I__1229\ : IoSpan4Mux
    port map (
            O => \N__5643\,
            I => \N__5637\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__5640\,
            I => \A_c_29\
        );

    \I__1227\ : Odrv4
    port map (
            O => \N__5637\,
            I => \A_c_29\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5628\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5631\,
            I => \N__5624\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5628\,
            I => \N__5621\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5627\,
            I => \N__5618\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5624\,
            I => \N__5615\
        );

    \I__1221\ : Span4Mux_v
    port map (
            O => \N__5621\,
            I => \N__5610\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5610\
        );

    \I__1219\ : Span12Mux_s8_h
    port map (
            O => \N__5615\,
            I => \N__5607\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__5610\,
            I => \N__5604\
        );

    \I__1217\ : Odrv12
    port map (
            O => \N__5607\,
            I => \A_c_28\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__5604\,
            I => \A_c_28\
        );

    \I__1215\ : IoInMux
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__1213\ : Span4Mux_s3_h
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__1212\ : Odrv4
    port map (
            O => \N__5590\,
            I => \RAM_SPACEm_i\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__5587\,
            I => \N__5582\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__5586\,
            I => \N__5578\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__5585\,
            I => \N__5574\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5569\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5581\,
            I => \N__5569\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5566\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5577\,
            I => \N__5562\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5558\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5569\,
            I => \N__5553\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5566\,
            I => \N__5553\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5565\,
            I => \N__5548\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5548\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5545\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5558\,
            I => \N__5542\
        );

    \I__1197\ : Span4Mux_h
    port map (
            O => \N__5553\,
            I => \N__5535\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5535\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5545\,
            I => \N__5535\
        );

    \I__1194\ : Span12Mux_s6_v
    port map (
            O => \N__5542\,
            I => \N__5532\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__5535\,
            I => \N__5529\
        );

    \I__1192\ : Odrv12
    port map (
            O => \N__5532\,
            I => \SIZ_c_1\
        );

    \I__1191\ : Odrv4
    port map (
            O => \N__5529\,
            I => \SIZ_c_1\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5510\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5523\,
            I => \N__5510\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5510\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5503\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5503\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5519\,
            I => \N__5503\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5518\,
            I => \N__5498\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5517\,
            I => \N__5498\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5510\,
            I => \U400_SDRAM.N_303_0_i\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__5503\,
            I => \U400_SDRAM.N_303_0_i\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5498\,
            I => \U400_SDRAM.N_303_0_i\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5485\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5485\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5485\,
            I => \U400_SDRAM.SDRAM_CMD_5_sqmuxa\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5482\,
            I => \N__5479\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5476\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__1173\ : Odrv4
    port map (
            O => \N__5473\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_1\
        );

    \I__1172\ : CEMux
    port map (
            O => \N__5470\,
            I => \N__5466\
        );

    \I__1171\ : CEMux
    port map (
            O => \N__5469\,
            I => \N__5463\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5466\,
            I => \N__5460\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__5463\,
            I => \N__5457\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__5460\,
            I => \N__5454\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__5457\,
            I => \N__5451\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__5454\,
            I => \U400_SDRAM.SDRAM_COUNTERe_0_i\
        );

    \I__1165\ : Odrv4
    port map (
            O => \N__5451\,
            I => \U400_SDRAM.SDRAM_COUNTERe_0_i\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5441\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5436\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5436\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5441\,
            I => \U400_SDRAM.N_66\
        );

    \I__1160\ : LocalMux
    port map (
            O => \N__5436\,
            I => \U400_SDRAM.N_66\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5427\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5422\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__5427\,
            I => \N__5419\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5426\,
            I => \N__5416\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5425\,
            I => \N__5413\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5422\,
            I => \U400_SDRAM.N_55\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__5419\,
            I => \U400_SDRAM.N_55\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5416\,
            I => \U400_SDRAM.N_55\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5413\,
            I => \U400_SDRAM.N_55\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5404\,
            I => \N__5400\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5403\,
            I => \N__5397\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5400\,
            I => \N__5394\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5397\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__5394\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__5389\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5380\,
            I => \N__5377\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__5377\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0\
        );

    \I__1140\ : InMux
    port map (
            O => \N__5374\,
            I => \N__5367\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5360\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5360\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5360\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5370\,
            I => \N__5356\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5367\,
            I => \N__5353\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__5360\,
            I => \N__5350\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5347\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__5356\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__1131\ : Odrv4
    port map (
            O => \N__5353\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__5350\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__5347\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5338\,
            I => \N__5326\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5337\,
            I => \N__5321\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5336\,
            I => \N__5321\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5316\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5334\,
            I => \N__5316\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__5333\,
            I => \N__5311\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5305\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__5331\,
            I => \N__5300\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5295\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5329\,
            I => \N__5295\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5326\,
            I => \N__5292\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__5321\,
            I => \N__5287\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5316\,
            I => \N__5287\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5315\,
            I => \N__5282\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5282\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5279\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5276\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5271\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5271\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5305\,
            I => \N__5268\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5261\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5261\
        );

    \I__1106\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5261\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5295\,
            I => \N__5258\
        );

    \I__1104\ : Span4Mux_v
    port map (
            O => \N__5292\,
            I => \N__5251\
        );

    \I__1103\ : Span4Mux_v
    port map (
            O => \N__5287\,
            I => \N__5251\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5282\,
            I => \N__5251\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5279\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5276\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5271\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1098\ : Odrv4
    port map (
            O => \N__5268\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5261\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1096\ : Odrv4
    port map (
            O => \N__5258\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1095\ : Odrv4
    port map (
            O => \N__5251\,
            I => \U400_SDRAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__5236\,
            I => \N__5230\
        );

    \I__1093\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5224\
        );

    \I__1092\ : InMux
    port map (
            O => \N__5234\,
            I => \N__5217\
        );

    \I__1091\ : InMux
    port map (
            O => \N__5233\,
            I => \N__5217\
        );

    \I__1090\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5217\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5214\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__5228\,
            I => \N__5204\
        );

    \I__1087\ : InMux
    port map (
            O => \N__5227\,
            I => \N__5200\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5224\,
            I => \N__5193\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5193\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5193\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5213\,
            I => \N__5190\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5212\,
            I => \N__5186\
        );

    \I__1081\ : InMux
    port map (
            O => \N__5211\,
            I => \N__5183\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5176\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5176\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5171\
        );

    \I__1077\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5171\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5168\
        );

    \I__1075\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5165\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__5200\,
            I => \N__5161\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__5193\,
            I => \N__5156\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__5190\,
            I => \N__5156\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5153\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__5186\,
            I => \N__5148\
        );

    \I__1069\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5148\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5145\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5142\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5176\,
            I => \N__5135\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5171\,
            I => \N__5135\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5135\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5165\,
            I => \N__5132\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5164\,
            I => \N__5129\
        );

    \I__1061\ : Span4Mux_v
    port map (
            O => \N__5161\,
            I => \N__5126\
        );

    \I__1060\ : Span4Mux_v
    port map (
            O => \N__5156\,
            I => \N__5123\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5120\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__5148\,
            I => \N__5113\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5145\,
            I => \N__5113\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5142\,
            I => \N__5113\
        );

    \I__1055\ : Span4Mux_h
    port map (
            O => \N__5135\,
            I => \N__5106\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__5132\,
            I => \N__5106\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__5129\,
            I => \N__5106\
        );

    \I__1052\ : Span4Mux_h
    port map (
            O => \N__5126\,
            I => \N__5099\
        );

    \I__1051\ : Span4Mux_h
    port map (
            O => \N__5123\,
            I => \N__5099\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__5120\,
            I => \N__5099\
        );

    \I__1049\ : Span4Mux_v
    port map (
            O => \N__5113\,
            I => \N__5096\
        );

    \I__1048\ : Span4Mux_v
    port map (
            O => \N__5106\,
            I => \N__5093\
        );

    \I__1047\ : Span4Mux_h
    port map (
            O => \N__5099\,
            I => \N__5090\
        );

    \I__1046\ : Span4Mux_h
    port map (
            O => \N__5096\,
            I => \N__5087\
        );

    \I__1045\ : Span4Mux_h
    port map (
            O => \N__5093\,
            I => \N__5084\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__5090\,
            I => \RESETn_c\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__5087\,
            I => \RESETn_c\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__5084\,
            I => \RESETn_c\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5069\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5069\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__5075\,
            I => \N__5063\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5053\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5069\,
            I => \N__5050\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5047\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5044\
        );

    \I__1034\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5041\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5063\,
            I => \N__5036\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5031\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5031\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5060\,
            I => \N__5024\
        );

    \I__1029\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5024\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5024\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5021\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5056\,
            I => \N__5018\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5053\,
            I => \N__5007\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__5050\,
            I => \N__5007\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5007\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5044\,
            I => \N__5007\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5041\,
            I => \N__5007\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5004\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5001\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5036\,
            I => \N__4994\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__4994\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__4994\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5021\,
            I => \N__4991\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5018\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1013\ : Odrv4
    port map (
            O => \N__5007\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5004\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5001\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1010\ : Odrv4
    port map (
            O => \N__4994\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__4991\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1008\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4968\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4965\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4976\,
            I => \N__4958\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4953\
        );

    \I__1004\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4953\
        );

    \I__1003\ : InMux
    port map (
            O => \N__4973\,
            I => \N__4947\
        );

    \I__1002\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4947\
        );

    \I__1001\ : InMux
    port map (
            O => \N__4971\,
            I => \N__4941\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4936\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__4965\,
            I => \N__4936\
        );

    \I__998\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4929\
        );

    \I__997\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4929\
        );

    \I__996\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4929\
        );

    \I__995\ : CascadeMux
    port map (
            O => \N__4961\,
            I => \N__4926\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4958\,
            I => \N__4919\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4953\,
            I => \N__4919\
        );

    \I__992\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4914\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__4947\,
            I => \N__4911\
        );

    \I__990\ : InMux
    port map (
            O => \N__4946\,
            I => \N__4904\
        );

    \I__989\ : InMux
    port map (
            O => \N__4945\,
            I => \N__4904\
        );

    \I__988\ : InMux
    port map (
            O => \N__4944\,
            I => \N__4904\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__4941\,
            I => \N__4897\
        );

    \I__986\ : Span4Mux_h
    port map (
            O => \N__4936\,
            I => \N__4897\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__4929\,
            I => \N__4897\
        );

    \I__984\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4890\
        );

    \I__983\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4890\
        );

    \I__982\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4890\
        );

    \I__981\ : Span4Mux_v
    port map (
            O => \N__4919\,
            I => \N__4887\
        );

    \I__980\ : InMux
    port map (
            O => \N__4918\,
            I => \N__4882\
        );

    \I__979\ : InMux
    port map (
            O => \N__4917\,
            I => \N__4882\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4914\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__977\ : Odrv4
    port map (
            O => \N__4911\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4904\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__975\ : Odrv4
    port map (
            O => \N__4897\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__4890\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__4887\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4882\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__971\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4861\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__4866\,
            I => \N__4858\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__4865\,
            I => \N__4853\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__4864\,
            I => \N__4849\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__4861\,
            I => \N__4842\
        );

    \I__966\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4839\
        );

    \I__965\ : CascadeMux
    port map (
            O => \N__4857\,
            I => \N__4834\
        );

    \I__964\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4828\
        );

    \I__963\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4828\
        );

    \I__962\ : InMux
    port map (
            O => \N__4852\,
            I => \N__4825\
        );

    \I__961\ : InMux
    port map (
            O => \N__4849\,
            I => \N__4822\
        );

    \I__960\ : InMux
    port map (
            O => \N__4848\,
            I => \N__4819\
        );

    \I__959\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4814\
        );

    \I__958\ : InMux
    port map (
            O => \N__4846\,
            I => \N__4814\
        );

    \I__957\ : InMux
    port map (
            O => \N__4845\,
            I => \N__4811\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__4842\,
            I => \N__4805\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4839\,
            I => \N__4805\
        );

    \I__954\ : InMux
    port map (
            O => \N__4838\,
            I => \N__4802\
        );

    \I__953\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4799\
        );

    \I__952\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4793\
        );

    \I__951\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4793\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__4828\,
            I => \N__4785\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4825\,
            I => \N__4785\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4822\,
            I => \N__4778\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4819\,
            I => \N__4778\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4814\,
            I => \N__4778\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__4811\,
            I => \N__4775\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \N__4771\
        );

    \I__943\ : Span4Mux_v
    port map (
            O => \N__4805\,
            I => \N__4763\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4763\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__4799\,
            I => \N__4763\
        );

    \I__940\ : InMux
    port map (
            O => \N__4798\,
            I => \N__4760\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4793\,
            I => \N__4757\
        );

    \I__938\ : InMux
    port map (
            O => \N__4792\,
            I => \N__4750\
        );

    \I__937\ : InMux
    port map (
            O => \N__4791\,
            I => \N__4750\
        );

    \I__936\ : InMux
    port map (
            O => \N__4790\,
            I => \N__4750\
        );

    \I__935\ : Span4Mux_v
    port map (
            O => \N__4785\,
            I => \N__4743\
        );

    \I__934\ : Span4Mux_h
    port map (
            O => \N__4778\,
            I => \N__4743\
        );

    \I__933\ : Span4Mux_v
    port map (
            O => \N__4775\,
            I => \N__4743\
        );

    \I__932\ : InMux
    port map (
            O => \N__4774\,
            I => \N__4736\
        );

    \I__931\ : InMux
    port map (
            O => \N__4771\,
            I => \N__4736\
        );

    \I__930\ : InMux
    port map (
            O => \N__4770\,
            I => \N__4736\
        );

    \I__929\ : Span4Mux_h
    port map (
            O => \N__4763\,
            I => \N__4733\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__4760\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__4757\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__4750\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__4743\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__4736\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__4733\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4720\,
            I => \N__4708\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__4719\,
            I => \N__4705\
        );

    \I__920\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4702\
        );

    \I__919\ : InMux
    port map (
            O => \N__4717\,
            I => \N__4699\
        );

    \I__918\ : InMux
    port map (
            O => \N__4716\,
            I => \N__4694\
        );

    \I__917\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4694\
        );

    \I__916\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4688\
        );

    \I__915\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4684\
        );

    \I__914\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4681\
        );

    \I__913\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4674\
        );

    \I__912\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4674\
        );

    \I__911\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4674\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__4702\,
            I => \N__4665\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__4699\,
            I => \N__4665\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__4694\,
            I => \N__4665\
        );

    \I__907\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4660\
        );

    \I__906\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4660\
        );

    \I__905\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4657\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4688\,
            I => \N__4654\
        );

    \I__903\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4651\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4684\,
            I => \N__4648\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4643\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__4674\,
            I => \N__4640\
        );

    \I__899\ : InMux
    port map (
            O => \N__4673\,
            I => \N__4632\
        );

    \I__898\ : InMux
    port map (
            O => \N__4672\,
            I => \N__4632\
        );

    \I__897\ : Span4Mux_v
    port map (
            O => \N__4665\,
            I => \N__4627\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4660\,
            I => \N__4627\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4657\,
            I => \N__4618\
        );

    \I__894\ : Span4Mux_h
    port map (
            O => \N__4654\,
            I => \N__4618\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4618\
        );

    \I__892\ : Span4Mux_h
    port map (
            O => \N__4648\,
            I => \N__4618\
        );

    \I__891\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4613\
        );

    \I__890\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4613\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4643\,
            I => \N__4608\
        );

    \I__888\ : Span4Mux_h
    port map (
            O => \N__4640\,
            I => \N__4608\
        );

    \I__887\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4603\
        );

    \I__886\ : InMux
    port map (
            O => \N__4638\,
            I => \N__4603\
        );

    \I__885\ : InMux
    port map (
            O => \N__4637\,
            I => \N__4600\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__4632\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__4627\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__4618\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4613\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__880\ : Odrv4
    port map (
            O => \N__4608\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__4603\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__4600\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__877\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4582\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__874\ : InMux
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__4573\,
            I => \N__4569\
        );

    \I__872\ : InMux
    port map (
            O => \N__4572\,
            I => \N__4566\
        );

    \I__871\ : Span4Mux_h
    port map (
            O => \N__4569\,
            I => \N__4563\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4566\,
            I => \U400_SDRAM.N_299_2\
        );

    \I__869\ : Odrv4
    port map (
            O => \N__4563\,
            I => \U400_SDRAM.N_299_2\
        );

    \I__868\ : CascadeMux
    port map (
            O => \N__4558\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__4555\,
            I => \N__4550\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__4554\,
            I => \N__4547\
        );

    \I__865\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4543\
        );

    \I__864\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4536\
        );

    \I__863\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4536\
        );

    \I__862\ : InMux
    port map (
            O => \N__4546\,
            I => \N__4536\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4543\,
            I => \N__4533\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4536\,
            I => \N__4530\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__4533\,
            I => \U400_SDRAM.N_266_0\
        );

    \I__858\ : Odrv4
    port map (
            O => \N__4530\,
            I => \U400_SDRAM.N_266_0\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__4525\,
            I => \U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_\
        );

    \I__856\ : IoInMux
    port map (
            O => \N__4522\,
            I => \N__4519\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4519\,
            I => \N__4516\
        );

    \I__854\ : Span4Mux_s2_v
    port map (
            O => \N__4516\,
            I => \N__4513\
        );

    \I__853\ : Odrv4
    port map (
            O => \N__4513\,
            I => \U400_BYTE_ENABLE_un1_LLBEn_i\
        );

    \I__852\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4504\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__4504\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__4501\,
            I => \U400_SDRAM.N_321_0_cascade_\
        );

    \I__848\ : InMux
    port map (
            O => \N__4498\,
            I => \N__4495\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4495\,
            I => \U400_SDRAM.N_322_0\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \N__4485\
        );

    \I__845\ : InMux
    port map (
            O => \N__4491\,
            I => \N__4480\
        );

    \I__844\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4477\
        );

    \I__843\ : InMux
    port map (
            O => \N__4489\,
            I => \N__4474\
        );

    \I__842\ : InMux
    port map (
            O => \N__4488\,
            I => \N__4469\
        );

    \I__841\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4469\
        );

    \I__840\ : CascadeMux
    port map (
            O => \N__4484\,
            I => \N__4466\
        );

    \I__839\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4463\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4480\,
            I => \N__4460\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__4477\,
            I => \N__4453\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4474\,
            I => \N__4453\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4469\,
            I => \N__4453\
        );

    \I__834\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4450\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4463\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__832\ : Odrv4
    port map (
            O => \N__4460\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__4453\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4450\,
            I => \U400_SDRAM.WRITE_CYCLEZ0\
        );

    \I__829\ : InMux
    port map (
            O => \N__4441\,
            I => \N__4438\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4438\,
            I => \U400_SDRAM.N_320_0\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__826\ : InMux
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__4429\,
            I => \N__4426\
        );

    \I__824\ : Span4Mux_h
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__823\ : Odrv4
    port map (
            O => \N__4423\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_0\
        );

    \I__822\ : InMux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__4417\,
            I => \U400_SDRAM.N_88\
        );

    \I__820\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4411\,
            I => \N__4408\
        );

    \I__818\ : Span4Mux_h
    port map (
            O => \N__4408\,
            I => \N__4405\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__4405\,
            I => \U400_SDRAM.SDRAM_COUNTER_s_3\
        );

    \I__816\ : InMux
    port map (
            O => \N__4402\,
            I => \N__4399\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__814\ : Span4Mux_v
    port map (
            O => \N__4396\,
            I => \N__4393\
        );

    \I__813\ : Odrv4
    port map (
            O => \N__4393\,
            I => \U400_SDRAM.N_56\
        );

    \I__812\ : CascadeMux
    port map (
            O => \N__4390\,
            I => \U400_SDRAM.N_56_cascade_\
        );

    \I__811\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4383\
        );

    \I__810\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4383\,
            I => \U400_SDRAM.N_108\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4380\,
            I => \U400_SDRAM.N_108\
        );

    \I__807\ : CascadeMux
    port map (
            O => \N__4375\,
            I => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_\
        );

    \I__806\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4368\
        );

    \I__805\ : InMux
    port map (
            O => \N__4371\,
            I => \N__4362\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4368\,
            I => \N__4359\
        );

    \I__803\ : InMux
    port map (
            O => \N__4367\,
            I => \N__4354\
        );

    \I__802\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4354\
        );

    \I__801\ : InMux
    port map (
            O => \N__4365\,
            I => \N__4351\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4362\,
            I => \U400_SDRAM.N_94_1\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__4359\,
            I => \U400_SDRAM.N_94_1\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4354\,
            I => \U400_SDRAM.N_94_1\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__4351\,
            I => \U400_SDRAM.N_94_1\
        );

    \I__796\ : CascadeMux
    port map (
            O => \N__4342\,
            I => \U400_SDRAM.N_275_cascade_\
        );

    \I__795\ : InMux
    port map (
            O => \N__4339\,
            I => \N__4332\
        );

    \I__794\ : InMux
    port map (
            O => \N__4338\,
            I => \N__4332\
        );

    \I__793\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4323\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4332\,
            I => \N__4320\
        );

    \I__791\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4315\
        );

    \I__790\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4315\
        );

    \I__789\ : InMux
    port map (
            O => \N__4329\,
            I => \N__4312\
        );

    \I__788\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4307\
        );

    \I__787\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4307\
        );

    \I__786\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4304\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4323\,
            I => \U400_SDRAM.N_54\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__4320\,
            I => \U400_SDRAM.N_54\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4315\,
            I => \U400_SDRAM.N_54\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4312\,
            I => \U400_SDRAM.N_54\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4307\,
            I => \U400_SDRAM.N_54\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4304\,
            I => \U400_SDRAM.N_54\
        );

    \I__779\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4288\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4288\,
            I => \U400_SDRAM.N_276\
        );

    \I__777\ : InMux
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__775\ : Span4Mux_h
    port map (
            O => \N__4279\,
            I => \N__4276\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__773\ : Span4Mux_v
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__772\ : Odrv4
    port map (
            O => \N__4270\,
            I => \A_c_26\
        );

    \I__771\ : IoInMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__769\ : Odrv12
    port map (
            O => \N__4261\,
            I => \MA_c_12\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__767\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__765\ : Span12Mux_v
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__764\ : Odrv12
    port map (
            O => \N__4246\,
            I => \A_c_20\
        );

    \I__763\ : IoInMux
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4240\,
            I => \N__4237\
        );

    \I__761\ : Span4Mux_s3_v
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__4234\,
            I => \MA_c_10\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__758\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4225\,
            I => \U400_SDRAM.N_30_2\
        );

    \I__756\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4219\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1\
        );

    \I__754\ : CascadeMux
    port map (
            O => \N__4216\,
            I => \U400_SDRAM.SDRAM_COUNTER44_5_cascade_\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__4213\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_\
        );

    \I__752\ : InMux
    port map (
            O => \N__4210\,
            I => \N__4207\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__750\ : Odrv12
    port map (
            O => \N__4204\,
            I => \U400_SDRAM.N_117\
        );

    \I__749\ : CascadeMux
    port map (
            O => \N__4201\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__4198\,
            I => \N__4195\
        );

    \I__747\ : InMux
    port map (
            O => \N__4195\,
            I => \N__4192\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__745\ : Odrv12
    port map (
            O => \N__4189\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4\
        );

    \I__744\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4182\
        );

    \I__743\ : InMux
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4182\,
            I => \U400_SDRAM.SDRAM_COUNTER42\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4179\,
            I => \U400_SDRAM.SDRAM_COUNTER42\
        );

    \I__740\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4170\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__4173\,
            I => \N__4167\
        );

    \I__738\ : LocalMux
    port map (
            O => \N__4170\,
            I => \N__4164\
        );

    \I__737\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4161\
        );

    \I__736\ : Odrv4
    port map (
            O => \N__4164\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER44_0\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4161\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER44_0\
        );

    \I__734\ : InMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4153\,
            I => \U400_SDRAM.TACK_4_m\
        );

    \I__732\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__730\ : Odrv12
    port map (
            O => \N__4144\,
            I => \U400_SDRAM.TACK_7_0\
        );

    \I__729\ : InMux
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__727\ : Span4Mux_h
    port map (
            O => \N__4135\,
            I => \N__4130\
        );

    \I__726\ : InMux
    port map (
            O => \N__4134\,
            I => \N__4122\
        );

    \I__725\ : InMux
    port map (
            O => \N__4133\,
            I => \N__4122\
        );

    \I__724\ : Span4Mux_h
    port map (
            O => \N__4130\,
            I => \N__4119\
        );

    \I__723\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4116\
        );

    \I__722\ : InMux
    port map (
            O => \N__4128\,
            I => \N__4111\
        );

    \I__721\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4111\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4122\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__719\ : Odrv4
    port map (
            O => \N__4119\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__4116\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4111\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_2\
        );

    \I__716\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__714\ : Odrv12
    port map (
            O => \N__4096\,
            I => \U400_SDRAM.TA_EN11_m\
        );

    \I__713\ : InMux
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__4087\,
            I => \U400_SDRAM.un1_TA_COUNTER26_2_0\
        );

    \I__710\ : IoInMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__708\ : IoSpan4Mux
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__707\ : IoSpan4Mux
    port map (
            O => \N__4075\,
            I => \N__4071\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__4074\,
            I => \N__4068\
        );

    \I__705\ : Span4Mux_s3_v
    port map (
            O => \N__4071\,
            I => \N__4065\
        );

    \I__704\ : InMux
    port map (
            O => \N__4068\,
            I => \N__4062\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__4065\,
            I => \TA_OUT\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4062\,
            I => \TA_OUT\
        );

    \I__701\ : ClkMux
    port map (
            O => \N__4057\,
            I => \N__3961\
        );

    \I__700\ : ClkMux
    port map (
            O => \N__4056\,
            I => \N__3961\
        );

    \I__699\ : ClkMux
    port map (
            O => \N__4055\,
            I => \N__3961\
        );

    \I__698\ : ClkMux
    port map (
            O => \N__4054\,
            I => \N__3961\
        );

    \I__697\ : ClkMux
    port map (
            O => \N__4053\,
            I => \N__3961\
        );

    \I__696\ : ClkMux
    port map (
            O => \N__4052\,
            I => \N__3961\
        );

    \I__695\ : ClkMux
    port map (
            O => \N__4051\,
            I => \N__3961\
        );

    \I__694\ : ClkMux
    port map (
            O => \N__4050\,
            I => \N__3961\
        );

    \I__693\ : ClkMux
    port map (
            O => \N__4049\,
            I => \N__3961\
        );

    \I__692\ : ClkMux
    port map (
            O => \N__4048\,
            I => \N__3961\
        );

    \I__691\ : ClkMux
    port map (
            O => \N__4047\,
            I => \N__3961\
        );

    \I__690\ : ClkMux
    port map (
            O => \N__4046\,
            I => \N__3961\
        );

    \I__689\ : ClkMux
    port map (
            O => \N__4045\,
            I => \N__3961\
        );

    \I__688\ : ClkMux
    port map (
            O => \N__4044\,
            I => \N__3961\
        );

    \I__687\ : ClkMux
    port map (
            O => \N__4043\,
            I => \N__3961\
        );

    \I__686\ : ClkMux
    port map (
            O => \N__4042\,
            I => \N__3961\
        );

    \I__685\ : ClkMux
    port map (
            O => \N__4041\,
            I => \N__3961\
        );

    \I__684\ : ClkMux
    port map (
            O => \N__4040\,
            I => \N__3961\
        );

    \I__683\ : ClkMux
    port map (
            O => \N__4039\,
            I => \N__3961\
        );

    \I__682\ : ClkMux
    port map (
            O => \N__4038\,
            I => \N__3961\
        );

    \I__681\ : ClkMux
    port map (
            O => \N__4037\,
            I => \N__3961\
        );

    \I__680\ : ClkMux
    port map (
            O => \N__4036\,
            I => \N__3961\
        );

    \I__679\ : ClkMux
    port map (
            O => \N__4035\,
            I => \N__3961\
        );

    \I__678\ : ClkMux
    port map (
            O => \N__4034\,
            I => \N__3961\
        );

    \I__677\ : ClkMux
    port map (
            O => \N__4033\,
            I => \N__3961\
        );

    \I__676\ : ClkMux
    port map (
            O => \N__4032\,
            I => \N__3961\
        );

    \I__675\ : ClkMux
    port map (
            O => \N__4031\,
            I => \N__3961\
        );

    \I__674\ : ClkMux
    port map (
            O => \N__4030\,
            I => \N__3961\
        );

    \I__673\ : ClkMux
    port map (
            O => \N__4029\,
            I => \N__3961\
        );

    \I__672\ : ClkMux
    port map (
            O => \N__4028\,
            I => \N__3961\
        );

    \I__671\ : ClkMux
    port map (
            O => \N__4027\,
            I => \N__3961\
        );

    \I__670\ : ClkMux
    port map (
            O => \N__4026\,
            I => \N__3961\
        );

    \I__669\ : GlobalMux
    port map (
            O => \N__3961\,
            I => \N__3958\
        );

    \I__668\ : gio2CtrlBuf
    port map (
            O => \N__3958\,
            I => \CLK40_c_g\
        );

    \I__667\ : InMux
    port map (
            O => \N__3955\,
            I => \N__3951\
        );

    \I__666\ : InMux
    port map (
            O => \N__3954\,
            I => \N__3948\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__3951\,
            I => \N__3944\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3948\,
            I => \N__3939\
        );

    \I__663\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3934\
        );

    \I__662\ : Span4Mux_v
    port map (
            O => \N__3944\,
            I => \N__3931\
        );

    \I__661\ : InMux
    port map (
            O => \N__3943\,
            I => \N__3926\
        );

    \I__660\ : InMux
    port map (
            O => \N__3942\,
            I => \N__3926\
        );

    \I__659\ : Span4Mux_h
    port map (
            O => \N__3939\,
            I => \N__3923\
        );

    \I__658\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3920\
        );

    \I__657\ : InMux
    port map (
            O => \N__3937\,
            I => \N__3917\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__3934\,
            I => \U400_SDRAM.N_105\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__3931\,
            I => \U400_SDRAM.N_105\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3926\,
            I => \U400_SDRAM.N_105\
        );

    \I__653\ : Odrv4
    port map (
            O => \N__3923\,
            I => \U400_SDRAM.N_105\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__3920\,
            I => \U400_SDRAM.N_105\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3917\,
            I => \U400_SDRAM.N_105\
        );

    \I__650\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3900\
        );

    \I__649\ : InMux
    port map (
            O => \N__3903\,
            I => \N__3897\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3900\,
            I => \N__3892\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3897\,
            I => \N__3889\
        );

    \I__646\ : InMux
    port map (
            O => \N__3896\,
            I => \N__3886\
        );

    \I__645\ : InMux
    port map (
            O => \N__3895\,
            I => \N__3883\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__3892\,
            I => \U400_SDRAM.N_59\
        );

    \I__643\ : Odrv12
    port map (
            O => \N__3889\,
            I => \U400_SDRAM.N_59\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3886\,
            I => \U400_SDRAM.N_59\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3883\,
            I => \U400_SDRAM.N_59\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3874\,
            I => \U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_\
        );

    \I__639\ : InMux
    port map (
            O => \N__3871\,
            I => \N__3868\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3868\,
            I => \U400_SDRAM.N_84\
        );

    \I__637\ : InMux
    port map (
            O => \N__3865\,
            I => \N__3861\
        );

    \I__636\ : InMux
    port map (
            O => \N__3864\,
            I => \N__3858\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3861\,
            I => \N__3855\
        );

    \I__634\ : LocalMux
    port map (
            O => \N__3858\,
            I => \N__3852\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__3855\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3852\,
            I => \U400_SDRAM.RAM_CYCLEZ0\
        );

    \I__631\ : CascadeMux
    port map (
            O => \N__3847\,
            I => \U400_SDRAM.N_30_2_cascade_\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__3844\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_\
        );

    \I__629\ : InMux
    port map (
            O => \N__3841\,
            I => \N__3838\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__3835\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0\
        );

    \I__626\ : InMux
    port map (
            O => \N__3832\,
            I => \N__3828\
        );

    \I__625\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3825\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3828\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3825\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__622\ : InMux
    port map (
            O => \N__3820\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\
        );

    \I__621\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3813\
        );

    \I__620\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3810\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3813\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3810\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__617\ : InMux
    port map (
            O => \N__3805\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\
        );

    \I__616\ : InMux
    port map (
            O => \N__3802\,
            I => \N__3798\
        );

    \I__615\ : InMux
    port map (
            O => \N__3801\,
            I => \N__3795\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3798\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3795\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__612\ : InMux
    port map (
            O => \N__3790\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\
        );

    \I__611\ : InMux
    port map (
            O => \N__3787\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\
        );

    \I__610\ : SRMux
    port map (
            O => \N__3784\,
            I => \N__3780\
        );

    \I__609\ : SRMux
    port map (
            O => \N__3783\,
            I => \N__3777\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3780\,
            I => \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3777\,
            I => \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\
        );

    \I__606\ : InMux
    port map (
            O => \N__3772\,
            I => \N__3769\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__3769\,
            I => \N__3766\
        );

    \I__604\ : Sp12to4
    port map (
            O => \N__3766\,
            I => \N__3763\
        );

    \I__603\ : Span12Mux_v
    port map (
            O => \N__3763\,
            I => \N__3760\
        );

    \I__602\ : Odrv12
    port map (
            O => \N__3760\,
            I => \A_c_24\
        );

    \I__601\ : CascadeMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__600\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__598\ : Span4Mux_v
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__597\ : Span4Mux_h
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__595\ : Odrv4
    port map (
            O => \N__3739\,
            I => \A_c_18\
        );

    \I__594\ : IoInMux
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__3730\,
            I => \MA_c_8\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__590\ : InMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__588\ : Sp12to4
    port map (
            O => \N__3718\,
            I => \N__3715\
        );

    \I__587\ : Span12Mux_s10_v
    port map (
            O => \N__3715\,
            I => \N__3712\
        );

    \I__586\ : Odrv12
    port map (
            O => \N__3712\,
            I => \A_c_19\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__3709\,
            I => \N__3706\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__3706\,
            I => \N__3703\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__3703\,
            I => \MA_c_9\
        );

    \I__582\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3697\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3697\,
            I => \N__3693\
        );

    \I__580\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3690\
        );

    \I__579\ : Span4Mux_v
    port map (
            O => \N__3693\,
            I => \N__3687\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3690\,
            I => \N__3684\
        );

    \I__577\ : Odrv4
    port map (
            O => \N__3687\,
            I => \U400_SDRAM.N_110\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__3684\,
            I => \U400_SDRAM.N_110\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__574\ : InMux
    port map (
            O => \N__3676\,
            I => \N__3673\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__572\ : Odrv12
    port map (
            O => \N__3670\,
            I => \RnW_c\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__570\ : InMux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3661\,
            I => \U400_SDRAM.N_57\
        );

    \I__568\ : InMux
    port map (
            O => \N__3658\,
            I => \N__3652\
        );

    \I__567\ : InMux
    port map (
            O => \N__3657\,
            I => \N__3652\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__3652\,
            I => \U400_SDRAM.N_51\
        );

    \I__565\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3645\
        );

    \I__564\ : InMux
    port map (
            O => \N__3648\,
            I => \N__3642\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3645\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__3642\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__3637\,
            I => \N__3634\
        );

    \I__560\ : InMux
    port map (
            O => \N__3634\,
            I => \N__3629\
        );

    \I__559\ : InMux
    port map (
            O => \N__3633\,
            I => \N__3624\
        );

    \I__558\ : InMux
    port map (
            O => \N__3632\,
            I => \N__3624\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3629\,
            I => \N__3621\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3624\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__555\ : Odrv4
    port map (
            O => \N__3621\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\
        );

    \I__554\ : InMux
    port map (
            O => \N__3616\,
            I => \N__3613\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__3613\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__552\ : InMux
    port map (
            O => \N__3610\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\
        );

    \I__551\ : InMux
    port map (
            O => \N__3607\,
            I => \N__3603\
        );

    \I__550\ : InMux
    port map (
            O => \N__3606\,
            I => \N__3600\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3603\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3600\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__547\ : InMux
    port map (
            O => \N__3595\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\
        );

    \I__546\ : InMux
    port map (
            O => \N__3592\,
            I => \N__3588\
        );

    \I__545\ : InMux
    port map (
            O => \N__3591\,
            I => \N__3585\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3588\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3585\,
            I => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__542\ : InMux
    port map (
            O => \N__3580\,
            I => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\
        );

    \I__541\ : InMux
    port map (
            O => \N__3577\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_6\
        );

    \I__540\ : InMux
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3571\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1\
        );

    \I__538\ : InMux
    port map (
            O => \N__3568\,
            I => \N__3562\
        );

    \I__537\ : InMux
    port map (
            O => \N__3567\,
            I => \N__3562\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3562\,
            I => \U400_SDRAM.N_111\
        );

    \I__535\ : InMux
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3556\,
            I => \N__3553\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__3553\,
            I => \N__3550\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3547\,
            I => \TSn_c\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3544\,
            I => \U400_SDRAM.un3_RAM_CYCLE_START_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3535\
        );

    \I__528\ : InMux
    port map (
            O => \N__3540\,
            I => \N__3535\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__526\ : Span4Mux_h
    port map (
            O => \N__3532\,
            I => \N__3523\
        );

    \I__525\ : InMux
    port map (
            O => \N__3531\,
            I => \N__3520\
        );

    \I__524\ : InMux
    port map (
            O => \N__3530\,
            I => \N__3517\
        );

    \I__523\ : InMux
    port map (
            O => \N__3529\,
            I => \N__3508\
        );

    \I__522\ : InMux
    port map (
            O => \N__3528\,
            I => \N__3508\
        );

    \I__521\ : InMux
    port map (
            O => \N__3527\,
            I => \N__3508\
        );

    \I__520\ : InMux
    port map (
            O => \N__3526\,
            I => \N__3508\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__3523\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3520\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3517\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3508\,
            I => \U400_SDRAM.RAM_CYCLE_STARTZ0\
        );

    \I__515\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3494\
        );

    \I__514\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3491\
        );

    \I__513\ : InMux
    port map (
            O => \N__3497\,
            I => \N__3488\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3494\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3491\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3488\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__509\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3476\
        );

    \I__508\ : InMux
    port map (
            O => \N__3480\,
            I => \N__3471\
        );

    \I__507\ : InMux
    port map (
            O => \N__3479\,
            I => \N__3471\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3476\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3471\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3466\,
            I => \N__3461\
        );

    \I__503\ : InMux
    port map (
            O => \N__3465\,
            I => \N__3458\
        );

    \I__502\ : InMux
    port map (
            O => \N__3464\,
            I => \N__3455\
        );

    \I__501\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3452\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3458\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3455\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3452\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__497\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3440\
        );

    \I__496\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3435\
        );

    \I__495\ : InMux
    port map (
            O => \N__3443\,
            I => \N__3435\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3440\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__3435\,
            I => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__492\ : CascadeMux
    port map (
            O => \N__3430\,
            I => \U400_SDRAM.N_54_cascade_\
        );

    \I__491\ : InMux
    port map (
            O => \N__3427\,
            I => \N__3424\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__3424\,
            I => \N__3421\
        );

    \I__489\ : Span12Mux_s11_h
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__488\ : Odrv12
    port map (
            O => \N__3418\,
            I => \A_c_9\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__3415\,
            I => \N__3412\
        );

    \I__486\ : InMux
    port map (
            O => \N__3412\,
            I => \N__3409\
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3409\,
            I => \N__3406\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__3406\,
            I => \N__3403\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3403\,
            I => \A_c_17\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__3400\,
            I => \N__3397\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3397\,
            I => \N__3394\
        );

    \I__480\ : Odrv12
    port map (
            O => \N__3394\,
            I => \MA_c_7\
        );

    \I__479\ : InMux
    port map (
            O => \N__3391\,
            I => \N__3388\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3388\,
            I => \N__3385\
        );

    \I__477\ : Odrv12
    port map (
            O => \N__3385\,
            I => \A_c_8\
        );

    \I__476\ : CascadeMux
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__475\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__472\ : Span4Mux_v
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3367\,
            I => \A_c_16\
        );

    \I__470\ : IoInMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3361\,
            I => \N__3358\
        );

    \I__468\ : Odrv12
    port map (
            O => \N__3358\,
            I => \MA_c_6\
        );

    \I__467\ : InMux
    port map (
            O => \N__3355\,
            I => \bfn_5_4_0_\
        );

    \I__466\ : InMux
    port map (
            O => \N__3352\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_0\
        );

    \I__465\ : InMux
    port map (
            O => \N__3349\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_1\
        );

    \I__464\ : InMux
    port map (
            O => \N__3346\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_2\
        );

    \I__463\ : InMux
    port map (
            O => \N__3343\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_3\
        );

    \I__462\ : InMux
    port map (
            O => \N__3340\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_4\
        );

    \I__461\ : InMux
    port map (
            O => \N__3337\,
            I => \U400_SDRAM.SDRAM_COUNTER_cry_5\
        );

    \I__460\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \U400_SDRAM.N_57_cascade_\
        );

    \I__459\ : InMux
    port map (
            O => \N__3331\,
            I => \N__3325\
        );

    \I__458\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3325\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3325\,
            I => \U400_SDRAM.N_46\
        );

    \I__456\ : CascadeMux
    port map (
            O => \N__3322\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_\
        );

    \I__455\ : CascadeMux
    port map (
            O => \N__3319\,
            I => \U400_SDRAM.N_266_0_cascade_\
        );

    \I__454\ : InMux
    port map (
            O => \N__3316\,
            I => \N__3312\
        );

    \I__453\ : InMux
    port map (
            O => \N__3315\,
            I => \N__3309\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3312\,
            I => \N__3303\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__3309\,
            I => \N__3303\
        );

    \I__450\ : InMux
    port map (
            O => \N__3308\,
            I => \N__3300\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__3303\,
            I => \U400_SDRAM.SDRAM_CMD12\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3300\,
            I => \U400_SDRAM.SDRAM_CMD12\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3295\,
            I => \U400_SDRAM.SDRAM_CMD12_cascade_\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__445\ : InMux
    port map (
            O => \N__3289\,
            I => \N__3283\
        );

    \I__444\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3283\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__3283\,
            I => \N__3280\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__3280\,
            I => \U400_SDRAM.un1_SDRAM_COUNTER52_0\
        );

    \I__441\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3273\
        );

    \I__440\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3270\
        );

    \I__439\ : LocalMux
    port map (
            O => \N__3273\,
            I => \N__3267\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3270\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__3267\,
            I => \U400_SDRAM.CS0_ENZ0\
        );

    \I__436\ : IoInMux
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3259\,
            I => \N__3256\
        );

    \I__434\ : IoSpan4Mux
    port map (
            O => \N__3256\,
            I => \N__3253\
        );

    \I__433\ : Span4Mux_s3_h
    port map (
            O => \N__3253\,
            I => \N__3250\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__3250\,
            I => \CS0n_c\
        );

    \I__431\ : IoInMux
    port map (
            O => \N__3247\,
            I => \N__3244\
        );

    \I__430\ : LocalMux
    port map (
            O => \N__3244\,
            I => \N__3241\
        );

    \I__429\ : Odrv12
    port map (
            O => \N__3241\,
            I => \WEn_c\
        );

    \I__428\ : IoInMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__426\ : Odrv12
    port map (
            O => \N__3232\,
            I => \CASn_c\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__424\ : InMux
    port map (
            O => \N__3226\,
            I => \N__3222\
        );

    \I__423\ : InMux
    port map (
            O => \N__3225\,
            I => \N__3219\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__3222\,
            I => \N__3216\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3219\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__420\ : Odrv12
    port map (
            O => \N__3216\,
            I => \U400_SDRAM.CS1_ENZ0\
        );

    \I__419\ : IoInMux
    port map (
            O => \N__3211\,
            I => \N__3208\
        );

    \I__418\ : LocalMux
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__417\ : IoSpan4Mux
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__416\ : Span4Mux_s3_v
    port map (
            O => \N__3202\,
            I => \N__3199\
        );

    \I__415\ : Odrv4
    port map (
            O => \N__3199\,
            I => \CS1n_c\
        );

    \I__414\ : CascadeMux
    port map (
            O => \N__3196\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__3193\,
            I => \U400_SDRAM.N_55_cascade_\
        );

    \I__412\ : CascadeMux
    port map (
            O => \N__3190\,
            I => \U400_SDRAM.N_105_cascade_\
        );

    \I__411\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3183\
        );

    \I__410\ : InMux
    port map (
            O => \N__3186\,
            I => \N__3180\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3183\,
            I => \U400_SDRAM.N_68\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3180\,
            I => \U400_SDRAM.N_68\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__3175\,
            I => \U400_SDRAM.N_62_cascade_\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3172\,
            I => \U400_SDRAM.N_39_cascade_\
        );

    \I__405\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3166\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3166\,
            I => \U400_SDRAM.N_62\
        );

    \I__403\ : CascadeMux
    port map (
            O => \N__3163\,
            I => \N__3160\
        );

    \I__402\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3154\
        );

    \I__401\ : InMux
    port map (
            O => \N__3159\,
            I => \N__3154\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3154\,
            I => \N__3151\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__3151\,
            I => \N__3148\
        );

    \I__398\ : Span4Mux_v
    port map (
            O => \N__3148\,
            I => \N__3145\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__3145\,
            I => \A_c_23\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3142\,
            I => \U400_SDRAM.N_41_cascade_\
        );

    \I__395\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3136\,
            I => \U400_SDRAM.N_52\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__3133\,
            I => \U400_SDRAM.N_295_0_cascade_\
        );

    \I__392\ : CascadeMux
    port map (
            O => \N__3130\,
            I => \U400_SDRAM.N_300_cascade_\
        );

    \I__391\ : InMux
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3124\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0\
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__3121\,
            I => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3118\,
            I => \U400_SDRAM.N_110_cascade_\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__3115\,
            I => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_\
        );

    \I__386\ : InMux
    port map (
            O => \N__3112\,
            I => \N__3107\
        );

    \I__385\ : InMux
    port map (
            O => \N__3111\,
            I => \N__3102\
        );

    \I__384\ : InMux
    port map (
            O => \N__3110\,
            I => \N__3102\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3107\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3102\,
            I => \U400_SDRAM.BURSTZ0\
        );

    \I__381\ : InMux
    port map (
            O => \N__3097\,
            I => \N__3088\
        );

    \I__380\ : InMux
    port map (
            O => \N__3096\,
            I => \N__3088\
        );

    \I__379\ : InMux
    port map (
            O => \N__3095\,
            I => \N__3084\
        );

    \I__378\ : InMux
    port map (
            O => \N__3094\,
            I => \N__3081\
        );

    \I__377\ : InMux
    port map (
            O => \N__3093\,
            I => \N__3078\
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3088\,
            I => \N__3075\
        );

    \I__375\ : InMux
    port map (
            O => \N__3087\,
            I => \N__3072\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__3084\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3081\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3078\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__3075\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3072\,
            I => \U400_SDRAM.TACKZ0\
        );

    \I__369\ : InMux
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__3055\,
            I => \N__3052\
        );

    \I__366\ : Odrv4
    port map (
            O => \N__3052\,
            I => \A_c_22\
        );

    \I__365\ : IoInMux
    port map (
            O => \N__3049\,
            I => \N__3046\
        );

    \I__364\ : LocalMux
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__363\ : IoSpan4Mux
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__362\ : Span4Mux_s1_h
    port map (
            O => \N__3040\,
            I => \N__3036\
        );

    \I__361\ : InMux
    port map (
            O => \N__3039\,
            I => \N__3033\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3036\,
            I => \BANK1_c\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__3033\,
            I => \BANK1_c\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__3028\,
            I => \N__3025\
        );

    \I__357\ : InMux
    port map (
            O => \N__3025\,
            I => \N__3022\
        );

    \I__356\ : LocalMux
    port map (
            O => \N__3022\,
            I => \N__3019\
        );

    \I__355\ : Span4Mux_v
    port map (
            O => \N__3019\,
            I => \N__3016\
        );

    \I__354\ : Odrv4
    port map (
            O => \N__3016\,
            I => \A_c_21\
        );

    \I__353\ : IoInMux
    port map (
            O => \N__3013\,
            I => \N__3010\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__351\ : Span12Mux_s1_h
    port map (
            O => \N__3007\,
            I => \N__3003\
        );

    \I__350\ : InMux
    port map (
            O => \N__3006\,
            I => \N__3000\
        );

    \I__349\ : Odrv12
    port map (
            O => \N__3003\,
            I => \BANK0_c\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3000\,
            I => \BANK0_c\
        );

    \I__347\ : IoInMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__345\ : Odrv4
    port map (
            O => \N__2989\,
            I => \RASn_c\
        );

    \I__344\ : CascadeMux
    port map (
            O => \N__2986\,
            I => \U400_SDRAM.N_299_cascade_\
        );

    \I__343\ : CascadeMux
    port map (
            O => \N__2983\,
            I => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__2980\,
            I => \U400_SDRAM.TA_COUNTER23_cascade_\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2977\,
            I => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2966\
        );

    \I__339\ : InMux
    port map (
            O => \N__2973\,
            I => \N__2963\
        );

    \I__338\ : InMux
    port map (
            O => \N__2972\,
            I => \N__2960\
        );

    \I__337\ : InMux
    port map (
            O => \N__2971\,
            I => \N__2953\
        );

    \I__336\ : InMux
    port map (
            O => \N__2970\,
            I => \N__2953\
        );

    \I__335\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2953\
        );

    \I__334\ : LocalMux
    port map (
            O => \N__2966\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__333\ : LocalMux
    port map (
            O => \N__2963\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__2960\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2953\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_1\
        );

    \I__330\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2932\
        );

    \I__329\ : InMux
    port map (
            O => \N__2943\,
            I => \N__2932\
        );

    \I__328\ : InMux
    port map (
            O => \N__2942\,
            I => \N__2929\
        );

    \I__327\ : InMux
    port map (
            O => \N__2941\,
            I => \N__2918\
        );

    \I__326\ : InMux
    port map (
            O => \N__2940\,
            I => \N__2918\
        );

    \I__325\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2918\
        );

    \I__324\ : InMux
    port map (
            O => \N__2938\,
            I => \N__2918\
        );

    \I__323\ : InMux
    port map (
            O => \N__2937\,
            I => \N__2918\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2932\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__321\ : LocalMux
    port map (
            O => \N__2929\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2918\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_0\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__2911\,
            I => \N__2905\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__2910\,
            I => \N__2901\
        );

    \I__317\ : CascadeMux
    port map (
            O => \N__2909\,
            I => \N__2898\
        );

    \I__316\ : CascadeMux
    port map (
            O => \N__2908\,
            I => \N__2895\
        );

    \I__315\ : InMux
    port map (
            O => \N__2905\,
            I => \N__2892\
        );

    \I__314\ : InMux
    port map (
            O => \N__2904\,
            I => \N__2889\
        );

    \I__313\ : InMux
    port map (
            O => \N__2901\,
            I => \N__2886\
        );

    \I__312\ : InMux
    port map (
            O => \N__2898\,
            I => \N__2881\
        );

    \I__311\ : InMux
    port map (
            O => \N__2895\,
            I => \N__2881\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2892\,
            I => \N__2878\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__2889\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2886\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2881\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__306\ : Odrv4
    port map (
            O => \N__2878\,
            I => \U400_SDRAM.TA_COUNTERZ0Z_3\
        );

    \I__305\ : InMux
    port map (
            O => \N__2869\,
            I => \N__2865\
        );

    \I__304\ : InMux
    port map (
            O => \N__2868\,
            I => \N__2862\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2865\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2862\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa\
        );

    \I__301\ : InMux
    port map (
            O => \N__2857\,
            I => \N__2853\
        );

    \I__300\ : CascadeMux
    port map (
            O => \N__2856\,
            I => \N__2850\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2853\,
            I => \N__2845\
        );

    \I__298\ : InMux
    port map (
            O => \N__2850\,
            I => \N__2842\
        );

    \I__297\ : InMux
    port map (
            O => \N__2849\,
            I => \N__2839\
        );

    \I__296\ : InMux
    port map (
            O => \N__2848\,
            I => \N__2836\
        );

    \I__295\ : Odrv4
    port map (
            O => \N__2845\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2842\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__293\ : LocalMux
    port map (
            O => \N__2839\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2836\,
            I => \U400_SDRAM.TA_COUNTER23\
        );

    \I__291\ : InMux
    port map (
            O => \N__2827\,
            I => \N__2823\
        );

    \I__290\ : InMux
    port map (
            O => \N__2826\,
            I => \N__2820\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2823\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2820\,
            I => \U400_SDRAM.TA_COUNTER27\
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2815\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\
        );

    \I__286\ : InMux
    port map (
            O => \N__2812\,
            I => \N__2809\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2809\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\
        );

    \I__284\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2803\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2803\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\
        );

    \I__282\ : CascadeMux
    port map (
            O => \N__2800\,
            I => \N__2797\
        );

    \I__281\ : InMux
    port map (
            O => \N__2797\,
            I => \N__2791\
        );

    \I__280\ : InMux
    port map (
            O => \N__2796\,
            I => \N__2791\
        );

    \I__279\ : LocalMux
    port map (
            O => \N__2791\,
            I => \U400_SDRAM.CO1\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2788\,
            I => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\
        );

    \I__277\ : CEMux
    port map (
            O => \N__2785\,
            I => \N__2782\
        );

    \I__276\ : LocalMux
    port map (
            O => \N__2782\,
            I => \N__2779\
        );

    \I__275\ : Span4Mux_s1_h
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__274\ : Odrv4
    port map (
            O => \N__2776\,
            I => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\
        );

    \I__273\ : IoInMux
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2770\,
            I => \RESETn_c_i\
        );

    \I__271\ : IoInMux
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2764\,
            I => \CONSTANT_ONE_NET\
        );

    \I__269\ : InMux
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__267\ : Odrv4
    port map (
            O => \N__2755\,
            I => \A_c_31\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__265\ : InMux
    port map (
            O => \N__2749\,
            I => \N__2746\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2746\,
            I => \N__2743\
        );

    \I__263\ : Span4Mux_h
    port map (
            O => \N__2743\,
            I => \N__2740\
        );

    \I__262\ : Odrv4
    port map (
            O => \N__2740\,
            I => \A_c_30\
        );

    \I__261\ : InMux
    port map (
            O => \N__2737\,
            I => \N__2734\
        );

    \I__260\ : LocalMux
    port map (
            O => \N__2734\,
            I => \N__2731\
        );

    \I__259\ : Odrv12
    port map (
            O => \N__2731\,
            I => \A_c_27\
        );

    \I__258\ : IoInMux
    port map (
            O => \N__2728\,
            I => \N__2725\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2725\,
            I => \N__2722\
        );

    \I__256\ : IoSpan4Mux
    port map (
            O => \N__2722\,
            I => \N__2719\
        );

    \I__255\ : Span4Mux_s3_h
    port map (
            O => \N__2719\,
            I => \N__2716\
        );

    \I__254\ : Span4Mux_h
    port map (
            O => \N__2716\,
            I => \N__2713\
        );

    \I__253\ : Span4Mux_h
    port map (
            O => \N__2713\,
            I => \N__2710\
        );

    \I__252\ : Span4Mux_v
    port map (
            O => \N__2710\,
            I => \N__2707\
        );

    \I__251\ : Odrv4
    port map (
            O => \N__2707\,
            I => \CLK40_ibuf_gb_io_gb_input\
        );

    \INVU400_SDRAM.MA_nesr_4C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_4C_net\,
            I => \N__4057\
        );

    \INVU400_SDRAM.MA_nesr_3C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_3C_net\,
            I => \N__4055\
        );

    \INVU400_SDRAM.MA_nesr_5C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_5C_net\,
            I => \N__4056\
        );

    \INVU400_SDRAM.MA_nesr_11C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_11C_net\,
            I => \N__4052\
        );

    \INVU400_SDRAM.SDRAM_CMD_1C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            I => \N__4045\
        );

    \INVU400_SDRAM.SDRAM_CONFIGUREDC\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            I => \N__4050\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            I => \N__4053\
        );

    \INVU400_SDRAM.MA_nesr_10C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_10C_net\,
            I => \N__4048\
        );

    \INVU400_SDRAM.MA_nesr_12C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_12C_net\,
            I => \N__4044\
        );

    \INVU400_SDRAM.RAM_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.RAM_CYCLEC_net\,
            I => \N__4049\
        );

    \INVU400_SDRAM.WRITE_CYCLEC\ : INV
    port map (
            O => \INVU400_SDRAM.WRITE_CYCLEC_net\,
            I => \N__4054\
        );

    \INVU400_SDRAM.MA_nesr_9C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_9C_net\,
            I => \N__4046\
        );

    \INVU400_SDRAM.MA_nesr_8C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_8C_net\,
            I => \N__4039\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            I => \N__4037\
        );

    \INVU400_SDRAM.REFRESH_COUNTER_0C\ : INV
    port map (
            O => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            I => \N__4040\
        );

    \INVU400_SDRAM.SDRAM_COUNTER_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            I => \N__4047\
        );

    \INVU400_SDRAM.MA_nesr_6C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_6C_net\,
            I => \N__4041\
        );

    \INVU400_SDRAM.MA_nesr_7C\ : INV
    port map (
            O => \INVU400_SDRAM.MA_nesr_7C_net\,
            I => \N__4035\
        );

    \INVU400_SDRAM.CS1nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS1nC_net\,
            I => \N__4032\
        );

    \INVU400_SDRAM.CS0nC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0nC_net\,
            I => \N__4027\
        );

    \INVU400_SDRAM.CS0_ENC\ : INV
    port map (
            O => \INVU400_SDRAM.CS0_ENC_net\,
            I => \N__4036\
        );

    \INVU400_SDRAM.SDRAM_CMD_0C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            I => \N__4038\
        );

    \INVU400_SDRAM.SDRAM_CMD_2C\ : INV
    port map (
            O => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            I => \N__4042\
        );

    \INVU400_SDRAM.RASnC\ : INV
    port map (
            O => \INVU400_SDRAM.RASnC_net\,
            I => \N__4026\
        );

    \INVU400_SDRAM.BANK1C\ : INV
    port map (
            O => \INVU400_SDRAM.BANK1C_net\,
            I => \N__4029\
        );

    \INVU400_SDRAM.TACKC\ : INV
    port map (
            O => \INVU400_SDRAM.TACKC_net\,
            I => \N__4031\
        );

    \INVU400_SDRAM.BURSTC\ : INV
    port map (
            O => \INVU400_SDRAM.BURSTC_net\,
            I => \N__4033\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_5_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_4_0_\
        );

    \CLK40_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2728\,
            GLOBALBUFFEROUTPUT => \CLK40_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2773\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_0_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6513\,
            in2 => \_gnd_net_\,
            in3 => \N__2812\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_1_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000000000000"
        )
    port map (
            in0 => \N__2974\,
            in1 => \N__2944\,
            in2 => \N__5236\,
            in3 => \N__2806\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_3_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110010000000"
        )
    port map (
            in0 => \N__4134\,
            in1 => \N__5234\,
            in2 => \N__2800\,
            in3 => \N__2904\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIJ78O_1_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2973\,
            in2 => \_gnd_net_\,
            in3 => \N__2943\,
            lcout => \U400_SDRAM.CO1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNI0LUG4_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__3093\,
            in1 => \N__2827\,
            in2 => \N__2856\,
            in3 => \N__2868\,
            lcout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0\,
            ltout => \U400_SDRAM.un1_TA_COUNTER_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_2_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__5233\,
            in1 => \N__2796\,
            in2 => \N__2788\,
            in3 => \N__4133\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4030\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011111111111"
        )
    port map (
            in0 => \N__2857\,
            in1 => \N__5227\,
            in2 => \_gnd_net_\,
            in3 => \N__3094\,
            lcout => \TA_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4028\,
            ce => \N__2785\,
            sr => \N__6479\
        );

    \RESETn_ibuf_RNIM9SF_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5213\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_3_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5235\,
            in1 => \N__2761\,
            in2 => \N__2752\,
            in3 => \N__2737\,
            lcout => \U400_ADDRESS_DECODE_RAM_SPACE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_3_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__2969\,
            in1 => \N__4127\,
            in2 => \N__2908\,
            in3 => \N__2937\,
            lcout => \U400_SDRAM.TA_COUNTER27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_2_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110010"
        )
    port map (
            in0 => \N__2971\,
            in1 => \N__4128\,
            in2 => \N__2909\,
            in3 => \N__2939\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_TA_COUNTER26_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_1_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001111"
        )
    port map (
            in0 => \N__3097\,
            in1 => \_gnd_net_\,
            in2 => \N__2983\,
            in3 => \N__2849\,
            lcout => \U400_SDRAM.un1_TA_COUNTER26_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_RNO_0_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2940\,
            in2 => \_gnd_net_\,
            in3 => \N__3112\,
            lcout => \U400_SDRAM.TA_EN11_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNIAJGG1_0_3_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__2938\,
            in1 => \N__4129\,
            in2 => \N__2910\,
            in3 => \N__2970\,
            lcout => \U400_SDRAM.TA_COUNTER23\,
            ltout => \U400_SDRAM.TA_COUNTER23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_RNO_0_0_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2941\,
            in2 => \N__2980\,
            in3 => \N__3096\,
            lcout => OPEN,
            ltout => \U400_SDRAM.TA_COUNTER_7_f1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_COUNTER_0_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2869\,
            in2 => \N__2977\,
            in3 => \N__5229\,
            lcout => \U400_SDRAM.TA_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4034\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST_RNISKH51_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__2972\,
            in1 => \N__2942\,
            in2 => \N__2911\,
            in3 => \N__3110\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa\,
            ltout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_EN_i_ess_RNO_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__2848\,
            in1 => \N__2826\,
            in2 => \N__2815\,
            in3 => \N__3087\,
            lcout => \U400_SDRAM.TA_COUNTER_0_sqmuxa_1_1_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__3111\,
            in1 => \N__3696\,
            in2 => \N__6352\,
            in3 => \N__3903\,
            lcout => \U400_SDRAM.BURSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BURSTC_net\,
            ce => 'H',
            sr => \N__6486\
        );

    \U400_SDRAM.TACK_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101100000001"
        )
    port map (
            in0 => \N__4210\,
            in1 => \N__4150\,
            in2 => \N__4198\,
            in3 => \N__3095\,
            lcout => \U400_SDRAM.TACKZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.TACKC_net\,
            ce => 'H',
            sr => \N__6482\
        );

    \U400_SDRAM.BANK1_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__3541\,
            in1 => \N__3061\,
            in2 => \N__3292\,
            in3 => \N__3039\,
            lcout => \BANK1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK1C_net\,
            ce => 'H',
            sr => \N__6480\
        );

    \U400_SDRAM.BANK0_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__3006\,
            in1 => \N__3288\,
            in2 => \N__3028\,
            in3 => \N__3540\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.BANK1C_net\,
            ce => 'H',
            sr => \N__6480\
        );

    \U400_SDRAM.RASn_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6835\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RASnC_net\,
            ce => 'H',
            sr => \N__6481\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_2_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000000"
        )
    port map (
            in0 => \N__4402\,
            in1 => \N__3315\,
            in2 => \N__4579\,
            in3 => \N__3530\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_299_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_2_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__6753\,
            in1 => \N__3127\,
            in2 => \N__2986\,
            in3 => \N__5904\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_2C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_2_LC_4_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3464\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3498\,
            lcout => \U400_SDRAM.N_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_5_2_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011011010"
        )
    port map (
            in0 => \N__5068\,
            in1 => \N__4977\,
            in2 => \N__4866\,
            in3 => \N__4714\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_295_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_2_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__3574\,
            in1 => \N__3139\,
            in2 => \N__3133\,
            in3 => \N__5336\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_300_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_2_LC_4_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5337\,
            in1 => \N__5074\,
            in2 => \N__3130\,
            in3 => \N__4510\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIQQB91_2_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__4846\,
            in1 => \N__5040\,
            in2 => \_gnd_net_\,
            in3 => \N__4327\,
            lcout => \U400_SDRAM.N_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_0_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111110"
        )
    port map (
            in0 => \N__4973\,
            in1 => \N__5430\,
            in2 => \N__4864\,
            in3 => \N__5335\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_0_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__6122\,
            in1 => \N__5903\,
            in2 => \N__3121\,
            in3 => \N__3841\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITAGQ1_1_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4693\,
            in2 => \_gnd_net_\,
            in3 => \N__3938\,
            lcout => \U400_SDRAM.N_110\,
            ltout => \U400_SDRAM.N_110_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNIFGBJ4_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__5209\,
            in1 => \N__3316\,
            in2 => \N__3118\,
            in3 => \N__3531\,
            lcout => \U400_SDRAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI5LLK_3_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__4972\,
            in1 => \N__4847\,
            in2 => \_gnd_net_\,
            in3 => \N__4692\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_a4_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNITM402_3_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110101"
        )
    port map (
            in0 => \N__5210\,
            in1 => \_gnd_net_\,
            in2 => \N__3115\,
            in3 => \N__4328\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_1_i_0_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI0TRC3_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5334\,
            in2 => \N__3196\,
            in3 => \N__3187\,
            lcout => \U400_SDRAM.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIFAF21_2_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5057\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4326\,
            lcout => \U400_SDRAM.N_55\,
            ltout => \U400_SDRAM.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIHPJJ1_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__5314\,
            in1 => \N__4837\,
            in2 => \N__3193\,
            in3 => \N__4974\,
            lcout => \U400_SDRAM.N_105\,
            ltout => \U400_SDRAM.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI2J773_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__4975\,
            in1 => \N__5315\,
            in2 => \N__3190\,
            in3 => \N__3186\,
            lcout => \U400_SDRAM.N_62\,
            ltout => \U400_SDRAM.N_62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_RNO_0_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__3159\,
            in1 => \N__4718\,
            in2 => \N__3175\,
            in3 => \N__3567\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_39_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0_EN_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111110111011"
        )
    port map (
            in0 => \N__3276\,
            in1 => \N__3330\,
            in2 => \N__3172\,
            in3 => \N__3657\,
            lcout => \U400_SDRAM.CS0_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6489\
        );

    \U400_SDRAM.CS1_EN_RNO_0_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4717\,
            in1 => \N__3169\,
            in2 => \N__3163\,
            in3 => \N__3568\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_41_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS1_EN_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111110111011"
        )
    port map (
            in0 => \N__3225\,
            in1 => \N__3331\,
            in2 => \N__3142\,
            in3 => \N__3658\,
            lcout => \U400_SDRAM.CS1_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0_ENC_net\,
            ce => 'H',
            sr => \N__6489\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI8E8G1_3_LC_4_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4867\,
            in1 => \N__4976\,
            in2 => \_gnd_net_\,
            in3 => \N__5425\,
            lcout => \U400_SDRAM.N_57\,
            ltout => \U400_SDRAM.N_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIG9NQ3_LC_4_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110010"
        )
    port map (
            in0 => \N__5338\,
            in1 => \N__3308\,
            in2 => \N__3334\,
            in3 => \N__4716\,
            lcout => \U400_SDRAM.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIJ1DL_6_LC_4_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3801\,
            in2 => \_gnd_net_\,
            in3 => \N__3816\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_o5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNI8CGL1_3_LC_4_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110000"
        )
    port map (
            in0 => \N__3606\,
            in1 => \N__3831\,
            in2 => \N__3322\,
            in3 => \N__3591\,
            lcout => \U400_SDRAM.N_266_0\,
            ltout => \U400_SDRAM.N_266_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIJU602_8_LC_4_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3319\,
            in3 => \N__5359\,
            lcout => \U400_SDRAM.SDRAM_CMD12\,
            ltout => \U400_SDRAM.SDRAM_CMD12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIG9NQ3_1_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4715\,
            in2 => \N__3295\,
            in3 => \N__3947\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.CS0n_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__6770\,
            in1 => \N__6308\,
            in2 => \N__6187\,
            in3 => \N__3277\,
            lcout => \CS0n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0nC_net\,
            ce => 'H',
            sr => \N__6487\
        );

    \U400_SDRAM.WEn_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6163\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0nC_net\,
            ce => 'H',
            sr => \N__6487\
        );

    \U400_SDRAM.CASn_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6309\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS0nC_net\,
            ce => 'H',
            sr => \N__6487\
        );

    \U400_SDRAM.CS1n_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__6771\,
            in1 => \N__6292\,
            in2 => \N__3229\,
            in3 => \N__6170\,
            lcout => \CS1n_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.CS1nC_net\,
            ce => 'H',
            sr => \N__6488\
        );

    \U400_SDRAM.MA_nesr_7_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3427\,
            in1 => \N__6772\,
            in2 => \N__3415\,
            in3 => \N__6659\,
            lcout => \MA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_7C_net\,
            ce => \N__6580\,
            sr => \N__6490\
        );

    \U400_SDRAM.MA_nesr_6_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3391\,
            in1 => \N__6776\,
            in2 => \N__3382\,
            in3 => \N__6667\,
            lcout => \MA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_6C_net\,
            ce => \N__6581\,
            sr => \N__6494\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_2_0_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4845\,
            in2 => \_gnd_net_\,
            in3 => \N__3355\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_5_4_0_\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_1_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4713\,
            in2 => \_gnd_net_\,
            in3 => \N__3352\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_0\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_2_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5522\,
            in1 => \N__5067\,
            in2 => \_gnd_net_\,
            in3 => \N__3349\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_1\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5469\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_3_LC_5_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4978\,
            in2 => \_gnd_net_\,
            in3 => \N__3346\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_s_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_2\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_4_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5523\,
            in1 => \N__3481\,
            in2 => \_gnd_net_\,
            in3 => \N__3343\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_3\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5469\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_5_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5517\,
            in1 => \N__3465\,
            in2 => \_gnd_net_\,
            in3 => \N__3340\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_4\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5469\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_6_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__3499\,
            in2 => \_gnd_net_\,
            in3 => \N__3337\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.SDRAM_COUNTER_cry_5\,
            carryout => \U400_SDRAM.SDRAM_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5469\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_7_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5518\,
            in1 => \N__3445\,
            in2 => \_gnd_net_\,
            in3 => \N__3577\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_2C_net\,
            ce => \N__5469\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNISRU82_8_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__5371\,
            in1 => \N__4546\,
            in2 => \_gnd_net_\,
            in3 => \N__3526\,
            lcout => \U400_SDRAM.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_0_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100000000"
        )
    port map (
            in0 => \N__3528\,
            in1 => \N__5373\,
            in2 => \N__4555\,
            in3 => \N__4367\,
            lcout => \U400_SDRAM.N_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_6_2_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5208\,
            in1 => \N__3480\,
            in2 => \_gnd_net_\,
            in3 => \N__3444\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_RNIDLIS3_8_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__3527\,
            in1 => \N__5372\,
            in2 => \N__4554\,
            in3 => \N__3937\,
            lcout => \U400_SDRAM.N_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_RNO_0_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__3559\,
            in1 => \N__5670\,
            in2 => \N__5710\,
            in3 => \N__5631\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un3_RAM_CYCLE_START_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_START_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001000000000"
        )
    port map (
            in0 => \N__3529\,
            in1 => \N__3864\,
            in2 => \N__3544\,
            in3 => \N__5207\,
            lcout => \U400_SDRAM.RAM_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4043\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI2OIR_7_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3497\,
            in1 => \N__3479\,
            in2 => \N__3466\,
            in3 => \N__3443\,
            lcout => \U400_SDRAM.N_54\,
            ltout => \U400_SDRAM.N_54_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIKV4N1_2_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4848\,
            in1 => \N__5039\,
            in2 => \N__3430\,
            in3 => \N__4366\,
            lcout => \U400_SDRAM.SDRAM_COUNTER42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNI24955_1_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__5404\,
            in1 => \N__3942\,
            in2 => \N__3667\,
            in3 => \N__4711\,
            lcout => \U400_SDRAM.N_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_3_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__4838\,
            in1 => \N__5426\,
            in2 => \N__4719\,
            in3 => \N__4489\,
            lcout => \U400_SDRAM.TACK_4_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2_1_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110110011"
        )
    port map (
            in0 => \N__3943\,
            in1 => \N__5189\,
            in2 => \N__4720\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_RNIJKCA2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_0_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3632\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__3783\
        );

    \U400_SDRAM.REFRESH_COUNTER_1_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__3633\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3649\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__3783\
        );

    \U400_SDRAM.un3_REFRESH_COUNTER_cry_1_c_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3648\,
            in2 => \N__3637\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.REFRESH_COUNTER_2_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3616\,
            in2 => \_gnd_net_\,
            in3 => \N__3610\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_1\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_3_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3607\,
            in2 => \_gnd_net_\,
            in3 => \N__3595\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_2\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_4_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3592\,
            in2 => \_gnd_net_\,
            in3 => \N__3580\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_3\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_5_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3832\,
            in2 => \_gnd_net_\,
            in3 => \N__3820\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_4\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_6_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3817\,
            in2 => \_gnd_net_\,
            in3 => \N__3805\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_5\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_7_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3802\,
            in2 => \_gnd_net_\,
            in3 => \N__3790\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \U400_SDRAM.un3_REFRESH_COUNTER_cry_6\,
            carryout => \U400_SDRAM.un3_REFRESH_COUNTER_cry_7\,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.REFRESH_COUNTER_8_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5370\,
            in2 => \_gnd_net_\,
            in3 => \N__3787\,
            lcout => \U400_SDRAM.REFRESH_COUNTERZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.REFRESH_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__3784\
        );

    \U400_SDRAM.MA_nesr_8_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3772\,
            in1 => \N__6823\,
            in2 => \N__3757\,
            in3 => \N__6658\,
            lcout => \MA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_8C_net\,
            ce => \N__6554\,
            sr => \N__6491\
        );

    \U400_SDRAM.SDRAM_CMD_RNIMFKP_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011011110111"
        )
    port map (
            in0 => \N__6821\,
            in1 => \N__6307\,
            in2 => \N__6517\,
            in3 => \N__6171\,
            lcout => \U400_SDRAM.un1_MA20_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_9_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6822\,
            in1 => \N__6306\,
            in2 => \N__3727\,
            in3 => \N__6196\,
            lcout => \MA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_9C_net\,
            ce => \N__6579\,
            sr => \N__6500\
        );

    \U400_SDRAM.WRITE_CYCLE_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000101110"
        )
    port map (
            in0 => \N__4483\,
            in1 => \N__3700\,
            in2 => \N__3679\,
            in3 => \N__3904\,
            lcout => \U400_SDRAM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.WRITE_CYCLEC_net\,
            ce => 'H',
            sr => \N__6502\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_0_0_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6402\,
            in1 => \N__3954\,
            in2 => \N__5585\,
            in3 => \N__3895\,
            lcout => \U400_SDRAM.N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TA_OUT_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__4141\,
            in1 => \N__4102\,
            in2 => \N__4074\,
            in3 => \N__4093\,
            lcout => \TA_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4051\,
            ce => 'H',
            sr => \N__6496\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNI8O963_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5212\,
            in1 => \N__4498\,
            in2 => \_gnd_net_\,
            in3 => \N__4337\,
            lcout => \U400_SDRAM.N_303_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIFGBJ4_1_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4672\,
            in1 => \N__3955\,
            in2 => \N__5228\,
            in3 => \N__3896\,
            lcout => \U400_SDRAM.SDRAM_CMD_5_sqmuxa\,
            ltout => \U400_SDRAM.SDRAM_CMD_5_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011011000"
        )
    port map (
            in0 => \N__4222\,
            in1 => \N__3865\,
            in2 => \N__3874\,
            in3 => \N__3871\,
            lcout => \U400_SDRAM.RAM_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.RAM_CYCLEC_net\,
            ce => 'H',
            sr => \N__6492\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIQ4PD_3_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4917\,
            in2 => \_gnd_net_\,
            in3 => \N__4637\,
            lcout => \U400_SDRAM.N_94_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIOLQ51_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__5056\,
            in1 => \N__5308\,
            in2 => \_gnd_net_\,
            in3 => \N__4329\,
            lcout => \U400_SDRAM.N_30_2\,
            ltout => \U400_SDRAM.N_30_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_0_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__5203\,
            in1 => \N__4185\,
            in2 => \N__3847\,
            in3 => \N__4371\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_0_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__4174\,
            in1 => \N__4490\,
            in2 => \N__3844\,
            in3 => \N__5309\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_i_a2_i_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.RAM_CYCLE_RNO_1_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111100"
        )
    port map (
            in0 => \N__4918\,
            in1 => \N__4798\,
            in2 => \N__4231\,
            in3 => \N__4673\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIN1PD_0_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4770\,
            in2 => \_gnd_net_\,
            in3 => \N__4638\,
            lcout => \U400_SDRAM.N_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNII7IR_2_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4639\,
            in1 => \N__5058\,
            in2 => \N__4810\,
            in3 => \N__4944\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_COUNTER44_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIPKQB2_3_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001110"
        )
    port map (
            in0 => \N__4945\,
            in1 => \N__5444\,
            in2 => \N__4216\,
            in3 => \N__4330\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER44_0\,
            ltout => \U400_SDRAM.un1_SDRAM_COUNTER44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_0_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4213\,
            in3 => \N__4488\,
            lcout => \U400_SDRAM.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNIPAEV_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5059\,
            in1 => \N__4774\,
            in2 => \N__4492\,
            in3 => \N__4365\,
            lcout => \U400_SDRAM.N_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_4_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100101111"
        )
    port map (
            in0 => \N__5445\,
            in1 => \N__5060\,
            in2 => \N__5333\,
            in3 => \N__4946\,
            lcout => OPEN,
            ltout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_2_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4387\,
            in2 => \N__4201\,
            in3 => \N__4331\,
            lcout => \U400_SDRAM.un1_SDRAM_COUNTER52_4_i_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.TACK_RNO_1_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010110001"
        )
    port map (
            in0 => \N__4491\,
            in1 => \N__4186\,
            in2 => \N__4173\,
            in3 => \N__4156\,
            lcout => \U400_SDRAM.TACK_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNIP3PD_3_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4852\,
            in2 => \_gnd_net_\,
            in3 => \N__4962\,
            lcout => \U400_SDRAM.N_56\,
            ltout => \U400_SDRAM.N_56_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_4_0_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110001000"
        )
    port map (
            in0 => \N__4964\,
            in1 => \N__5062\,
            in2 => \N__4390\,
            in3 => \N__4712\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_o2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_3_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4386\,
            in2 => \N__4375\,
            in3 => \N__4338\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_2_1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5332\,
            in1 => \N__4856\,
            in2 => \N__5075\,
            in3 => \N__4372\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_275_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_0_1_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101000"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__4291\,
            in2 => \N__4342\,
            in3 => \N__4339\,
            lcout => \U400_SDRAM.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__5061\,
            in1 => \N__4963\,
            in2 => \N__4865\,
            in3 => \N__4687\,
            lcout => \U400_SDRAM.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_12_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6188\,
            in1 => \N__4285\,
            in2 => \N__6310\,
            in3 => \N__6834\,
            lcout => \MA_c_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_12C_net\,
            ce => \N__6597\,
            sr => \N__6495\
        );

    \U400_SDRAM.MA_nesr_10_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__6847\,
            in1 => \N__6305\,
            in2 => \N__4258\,
            in3 => \N__6195\,
            lcout => \MA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_10C_net\,
            ce => \N__6569\,
            sr => \N__6501\
        );

    \U400_ADDRESS_DECODE.RAM_SPACE_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__5627\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__5709\,
            lcout => \RAM_SPACEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un2_LLBEn_0_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010000111100"
        )
    port map (
            in0 => \N__5760\,
            in1 => \N__6403\,
            in2 => \N__5587\,
            in3 => \N__5803\,
            lcout => OPEN,
            ltout => \U400_BYTE_ENABLE.un2_LLBEn_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LLBEn_i_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111110101"
        )
    port map (
            in0 => \N__5839\,
            in1 => \N__5759\,
            in2 => \N__4525\,
            in3 => \N__5581\,
            lcout => \U400_BYTE_ENABLE_un1_LLBEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_3_2_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__4925\,
            in1 => \N__4792\,
            in2 => \_gnd_net_\,
            in3 => \N__5211\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_76_i_a4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIE01O_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110001111110"
        )
    port map (
            in0 => \N__4647\,
            in1 => \N__4791\,
            in2 => \N__4961\,
            in3 => \N__5329\,
            lcout => OPEN,
            ltout => \U400_SDRAM.N_321_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIGMQQ1_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111110000"
        )
    port map (
            in0 => \N__5330\,
            in1 => \N__4441\,
            in2 => \N__4501\,
            in3 => \N__5066\,
            lcout => \U400_SDRAM.N_322_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.WRITE_CYCLE_RNICOHO_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000010011"
        )
    port map (
            in0 => \N__4790\,
            in1 => \N__4924\,
            in2 => \N__4484\,
            in3 => \N__4646\,
            lcout => \U400_SDRAM.N_320_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_0_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001110010"
        )
    port map (
            in0 => \N__5519\,
            in1 => \N__5380\,
            in2 => \N__4435\,
            in3 => \N__4420\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__5470\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5491\,
            in1 => \N__4414\,
            in2 => \N__6348\,
            in3 => \N__5521\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__5470\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_1_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__5490\,
            in2 => \N__6347\,
            in3 => \N__5482\,
            lcout => \U400_SDRAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_COUNTER_0C_net\,
            ce => \N__5470\,
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5304\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5403\,
            lcout => \U400_SDRAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CONFIGUREDC_net\,
            ce => 'H',
            sr => \N__6493\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNITAGQ1_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__4952\,
            in2 => \N__5331\,
            in3 => \N__5431\,
            lcout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U400_SDRAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_COUNTER_RNO_1_0_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__5182\,
            in1 => \N__5303\,
            in2 => \N__5389\,
            in3 => \N__5386\,
            lcout => \U400_SDRAM.SDRAM_COUNTER_cnst_0_a2_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_5_1_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5374\,
            in1 => \N__4833\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_a5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CONFIGURED_RNIVK7J_LC_7_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5310\,
            in1 => \N__5164\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U400_SDRAM.N_299_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_4_1_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__5077\,
            in1 => \N__4971\,
            in2 => \N__4857\,
            in3 => \N__4691\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNO_1_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101110011"
        )
    port map (
            in0 => \N__4585\,
            in1 => \N__4572\,
            in2 => \N__4558\,
            in3 => \N__4553\,
            lcout => OPEN,
            ltout => \U400_SDRAM.SDRAM_CMD_cnst_0_0_33_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__6255\,
            in1 => \N__5923\,
            in2 => \N__5914\,
            in3 => \N__5911\,
            lcout => \U400_SDRAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.SDRAM_CMD_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_11_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6842\,
            in1 => \N__6301\,
            in2 => \N__5887\,
            in3 => \N__6194\,
            lcout => \MA_c_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_11C_net\,
            ce => \N__6588\,
            sr => \N__6503\
        );

    \U400_BYTE_ENABLE.un1_UMBEn_i_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111100110011"
        )
    port map (
            in0 => \N__5765\,
            in1 => \N__5841\,
            in2 => \N__5586\,
            in3 => \N__5728\,
            lcout => \U400_BYTE_ENABLE_un1_UMBEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_LMBEn_i_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010101110101"
        )
    port map (
            in0 => \N__5840\,
            in1 => \N__5764\,
            in2 => \N__5722\,
            in3 => \N__5804\,
            lcout => \U400_BYTE_ENABLE_un1_LMBEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un1_UUBEn_i_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101100110011"
        )
    port map (
            in0 => \N__5766\,
            in1 => \N__5842\,
            in2 => \N__5811\,
            in3 => \N__5721\,
            lcout => \U400_BYTE_ENABLE_un1_UUBEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.un2_UMBEn_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111000100"
        )
    port map (
            in0 => \N__5812\,
            in1 => \N__6401\,
            in2 => \N__5767\,
            in3 => \N__5565\,
            lcout => \U400_BYTE_ENABLE.un2_UMBEn_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_BYTE_ENABLE.LW_TRANS_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__6400\,
            in1 => \_gnd_net_\,
            in2 => \N__5577\,
            in3 => \_gnd_net_\,
            lcout => \U400_BYTE_ENABLE.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_ADDRESS_DECODE.RAM_SPACEm_i_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__5705\,
            in1 => \N__5671\,
            in2 => \_gnd_net_\,
            in3 => \N__5632\,
            lcout => \RAM_SPACEm_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.BURST8_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6388\,
            lcout => \U400_SDRAM.BURSTZ0Z8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.SDRAM_CMD_RNI06O9_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6839\,
            in1 => \N__6286\,
            in2 => \_gnd_net_\,
            in3 => \N__6197\,
            lcout => \U400_SDRAM.MA19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_5_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100101110"
        )
    port map (
            in0 => \N__6198\,
            in1 => \N__6841\,
            in2 => \N__6322\,
            in3 => \N__6288\,
            lcout => \U400_SDRAM.MA_5_iv_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_RNO_0_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001110"
        )
    port map (
            in0 => \N__6840\,
            in1 => \N__6287\,
            in2 => \N__6214\,
            in3 => \N__6199\,
            lcout => \U400_SDRAM.MA_5_iv_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U400_SDRAM.MA_nesr_5_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6094\,
            in1 => \N__6082\,
            in2 => \_gnd_net_\,
            in3 => \N__6648\,
            lcout => \MA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_5C_net\,
            ce => \N__6593\,
            sr => \N__6505\
        );

    \U400_SDRAM.MA_nesr_3_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6061\,
            in1 => \N__6843\,
            in2 => \N__6052\,
            in3 => \N__6638\,
            lcout => \MA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_3C_net\,
            ce => \N__6592\,
            sr => \N__6504\
        );

    \U400_SDRAM.MA_nesr_4_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6846\,
            in1 => \N__6019\,
            in2 => \N__6007\,
            in3 => \N__6666\,
            lcout => \MA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_4C_net\,
            ce => \N__6598\,
            sr => \N__6506\
        );

    \U400_SDRAM.MA_nesr_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__6664\,
            in1 => \N__5974\,
            in2 => \N__5962\,
            in3 => \N__6844\,
            lcout => \MA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_4C_net\,
            ce => \N__6598\,
            sr => \N__6506\
        );

    \U400_SDRAM.MA_nesr_1_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__5938\,
            in1 => \N__5929\,
            in2 => \_gnd_net_\,
            in3 => \N__6663\,
            lcout => \MA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_4C_net\,
            ce => \N__6598\,
            sr => \N__6506\
        );

    \U400_SDRAM.MA_nesr_2_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__6845\,
            in1 => \N__6691\,
            in2 => \N__6679\,
            in3 => \N__6665\,
            lcout => \MA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU400_SDRAM.MA_nesr_4C_net\,
            ce => \N__6598\,
            sr => \N__6506\
        );

    \TAn_obuft_RNO_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_474_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

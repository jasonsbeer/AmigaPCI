-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Apr 20 2025 10:01:18

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    CMA : out std_logic_vector(10 downto 0);
    DA : out std_logic_vector(2 downto 0);
    A : in std_logic_vector(20 downto 0);
    DBRn : in std_logic;
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11999\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11845\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11827\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11791\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11782\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11439\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10893\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10702\ : std_logic;
signal \N__10699\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10681\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10529\ : std_logic;
signal \N__10526\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10369\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10360\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9967\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9756\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9747\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9582\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9573\ : std_logic;
signal \N__9570\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9534\ : std_logic;
signal \N__9531\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9228\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9186\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9036\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8996\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8988\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8832\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8409\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8238\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8133\ : std_logic;
signal \N__8124\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8016\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__7998\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7812\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7731\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7719\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7656\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7194\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7169\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7137\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6845\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6639\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6588\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6444\ : std_logic;
signal \N__6441\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6333\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6151\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6126\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5982\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5728\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5712\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5574\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5568\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5490\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5412\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5355\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5229\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5223\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5199\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5150\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4957\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4848\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4822\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4676\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4512\ : std_logic;
signal \N__4509\ : std_logic;
signal \N__4506\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4381\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4221\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4167\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4120\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4114\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4089\ : std_logic;
signal \N__4086\ : std_logic;
signal \N__4083\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4054\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \REGSPACEn_c\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ1Z_2\ : std_logic;
signal \U712_REG_SM.N_456\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_6_0_a2_0_a2_1_0\ : std_logic;
signal \U712_CHIP_RAM.N_607_cascade_\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_484\ : std_logic;
signal \U712_CHIP_RAM.N_607\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_480_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.REGENn_e_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_0\ : std_logic;
signal \U712_REG_SM.START_RSTZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\ : std_logic;
signal \U712_REG_SM.N_349_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CLK_EN_e_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_432_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_406_cascade_\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.N_515_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_326_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_614\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.N_614_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_3_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_338_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\ : std_logic;
signal \U712_CHIP_RAM.N_430_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_429\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_402_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_3\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \A_c_14\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CYCLE_TERM.N_486_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_EN6_0\ : std_logic;
signal \U712_REG_SM.N_465_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un3_DMA_CYCLE_START\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.N_347_cascade_\ : std_logic;
signal \U712_REG_SM.N_464\ : std_logic;
signal \U712_REG_SM.N_330\ : std_logic;
signal \U712_REG_SM.N_330_cascade_\ : std_logic;
signal \bfn_9_15_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_CHIP_RAM.N_471\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \U712_CHIP_RAM.N_477_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0\ : std_logic;
signal \U712_CHIP_RAM.N_406\ : std_logic;
signal \U712_CHIP_RAM.N_430\ : std_logic;
signal \U712_CHIP_RAM.N_44\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_500\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\ : std_logic;
signal \U712_CHIP_RAM.N_515\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_504_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_508_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_508\ : std_logic;
signal \U712_CHIP_RAM.N_610\ : std_logic;
signal \U712_CHIP_RAM.N_608\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_361\ : std_logic;
signal \CPU_TACKm\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_350\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTc_0_0\ : std_logic;
signal \U712_REG_SM.N_348_cascade_\ : std_logic;
signal \U712_REG_SM.N_347\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_4\ : std_logic;
signal \U712_REG_SM.N_399_cascade_\ : std_logic;
signal \U712_REG_SM.WRITE_CYCLEZ0\ : std_logic;
signal \U712_REG_SM.N_212\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ0Z_3\ : std_logic;
signal \U712_REG_SM.N_458\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.N_447\ : std_logic;
signal \RASn_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8\ : std_logic;
signal \A_c_17\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_432\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_4_cascade_\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_327\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_433\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.N_499\ : std_logic;
signal \U712_CHIP_RAM.N_499_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_341\ : std_logic;
signal \U712_CHIP_RAM.N_507_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_438\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.N_440_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_439\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.BANK0_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_507\ : std_logic;
signal \U712_CHIP_RAM.N_504\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_48\ : std_logic;
signal \LATCH_CLK_c\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_BYTE_ENABLE.N_443_cascade_\ : std_logic;
signal \N_32_i\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.BANK0_RNOZ0Z_3\ : std_logic;
signal \U712_REG_SM.STATE_COUNTZ1Z_2\ : std_logic;
signal \U712_REG_SM.N_348\ : std_logic;
signal \U712_REG_SM.N_462_cascade_\ : std_logic;
signal \U712_REG_SM.N_399\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_446\ : std_logic;
signal \N_435\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \CASn_c\ : std_logic;
signal \U712_CHIP_RAM.N_340\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\ : std_logic;
signal \U712_CHIP_RAM.DBENn_8_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \U712_CHIP_RAM.N_382\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U712_CHIP_RAM.N_374\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\ : std_logic;
signal \U712_CHIP_RAM.N_337\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_441\ : std_logic;
signal \N_34_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_451_cascade_\ : std_logic;
signal \N_200_i\ : std_logic;
signal \CPU_CYCLEm\ : std_logic;
signal \U712_BYTE_ENABLE.N_323_i\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \U712_BYTE_ENABLE.N_453_cascade_\ : std_logic;
signal \N_202_i\ : std_logic;
signal \CLK40_PLL_i\ : std_logic;
signal \CLK40_PLL_i_i\ : std_logic;
signal \N_334\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \ASn_c\ : std_logic;
signal \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \N_353_i\ : std_logic;
signal \N_354_i\ : std_logic;
signal \N_84_i\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_1\ : std_logic;
signal \N_355_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \WEn_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \U712_CHIP_RAM.N_501\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\ : std_logic;
signal \DMA_CYCLEm\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A1_nesrC_net\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \RnW_c\ : std_logic;
signal \WRITE_CYCLEm\ : std_logic;
signal \N_405\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \REG_CYCLEm\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \DA_wire\ : std_logic_vector(2 downto 0);
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    TBIn <= \TBIn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    DA <= \DA_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    TCIn <= \TCIn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL_i\,
            REFERENCECLK => \N__4072\,
            RESETB => \N__7360\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11999\,
            DIN => \N__11998\,
            DOUT => \N__11997\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11999\,
            PADOUT => \N__11998\,
            PADIN => \N__11997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11990\,
            DIN => \N__11989\,
            DOUT => \N__11988\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11990\,
            PADOUT => \N__11989\,
            PADIN => \N__11988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11981\,
            DIN => \N__11980\,
            DOUT => \N__11979\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11981\,
            PADOUT => \N__11980\,
            PADIN => \N__11979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7345\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11972\,
            DIN => \N__11971\,
            DOUT => \N__11970\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11972\,
            PADOUT => \N__11971\,
            PADIN => \N__11970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10129\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11963\,
            DIN => \N__11962\,
            DOUT => \N__11961\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11963\,
            PADOUT => \N__11962\,
            PADIN => \N__11961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11954\,
            DIN => \N__11953\,
            DOUT => \N__11952\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11954\,
            PADOUT => \N__11953\,
            PADIN => \N__11952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11945\,
            DIN => \N__11944\,
            DOUT => \N__11943\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11945\,
            PADOUT => \N__11944\,
            PADIN => \N__11943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11936\,
            DIN => \N__11935\,
            DOUT => \N__11934\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11936\,
            PADOUT => \N__11935\,
            PADIN => \N__11934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11927\,
            DIN => \N__11926\,
            DOUT => \N__11925\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11927\,
            PADOUT => \N__11926\,
            PADIN => \N__11925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11918\,
            DIN => \N__11917\,
            DOUT => \N__11916\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11918\,
            PADOUT => \N__11917\,
            PADIN => \N__11916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11909\,
            DIN => \N__11908\,
            DOUT => \N__11907\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11909\,
            PADOUT => \N__11908\,
            PADIN => \N__11907\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7030\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11900\,
            DIN => \N__11899\,
            DOUT => \N__11898\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11900\,
            PADOUT => \N__11899\,
            PADIN => \N__11898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8605\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11891\,
            DIN => \N__11890\,
            DOUT => \N__11889\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11891\,
            PADOUT => \N__11890\,
            PADIN => \N__11889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11882\,
            DIN => \N__11881\,
            DOUT => \N__11880\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11882\,
            PADOUT => \N__11881\,
            PADIN => \N__11880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11873\,
            DIN => \N__11872\,
            DOUT => \N__11871\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11873\,
            PADOUT => \N__11872\,
            PADIN => \N__11871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \REGSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11864\,
            DIN => \N__11863\,
            DOUT => \N__11862\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11864\,
            PADOUT => \N__11863\,
            PADIN => \N__11862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11855\,
            DIN => \N__11854\,
            DOUT => \N__11853\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11855\,
            PADOUT => \N__11854\,
            PADIN => \N__11853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5179\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11846\,
            DIN => \N__11845\,
            DOUT => \N__11844\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11846\,
            PADOUT => \N__11845\,
            PADIN => \N__11844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11837\,
            DIN => \N__11836\,
            DOUT => \N__11835\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11837\,
            PADOUT => \N__11836\,
            PADIN => \N__11835\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11828\,
            DIN => \N__11827\,
            DOUT => \N__11826\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11828\,
            PADOUT => \N__11827\,
            PADIN => \N__11826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8095\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11819\,
            DIN => \N__11818\,
            DOUT => \N__11817\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11819\,
            PADOUT => \N__11818\,
            PADIN => \N__11817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11810\,
            DIN => \N__11809\,
            DOUT => \N__11808\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11810\,
            PADOUT => \N__11809\,
            PADIN => \N__11808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9850\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11801\,
            DIN => \N__11800\,
            DOUT => \N__11799\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11801\,
            PADOUT => \N__11800\,
            PADIN => \N__11799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11792\,
            DIN => \N__11791\,
            DOUT => \N__11790\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11792\,
            PADOUT => \N__11791\,
            PADIN => \N__11790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8638\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11783\,
            DIN => \N__11782\,
            DOUT => \N__11781\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11783\,
            PADOUT => \N__11782\,
            PADIN => \N__11781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4711\,
            DIN0 => OPEN,
            DOUT0 => \N__4629\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11774\,
            DIN => \N__11773\,
            DOUT => \N__11772\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11774\,
            PADOUT => \N__11773\,
            PADIN => \N__11772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11765\,
            DIN => \N__11764\,
            DOUT => \N__11763\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11765\,
            PADOUT => \N__11764\,
            PADIN => \N__11763\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11756\,
            DIN => \N__11755\,
            DOUT => \N__11754\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11756\,
            PADOUT => \N__11755\,
            PADIN => \N__11754\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11747\,
            DIN => \N__11746\,
            DOUT => \N__11745\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11747\,
            PADOUT => \N__11746\,
            PADIN => \N__11745\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11738\,
            DIN => \N__11737\,
            DOUT => \N__11736\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11738\,
            PADOUT => \N__11737\,
            PADIN => \N__11736\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11729\,
            DIN => \N__11728\,
            DOUT => \N__11727\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11729\,
            PADOUT => \N__11728\,
            PADIN => \N__11727\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7378\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11720\,
            DIN => \N__11719\,
            DOUT => \N__11718\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11720\,
            PADOUT => \N__11719\,
            PADIN => \N__11718\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11711\,
            DIN => \N__11710\,
            DOUT => \N__11709\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11711\,
            PADOUT => \N__11710\,
            PADIN => \N__11709\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11702\,
            DIN => \N__11701\,
            DOUT => \N__11700\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11702\,
            PADOUT => \N__11701\,
            PADIN => \N__11700\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11693\,
            DIN => \N__11692\,
            DOUT => \N__11691\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11693\,
            PADOUT => \N__11692\,
            PADIN => \N__11691\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11684\,
            DIN => \N__11683\,
            DOUT => \N__11682\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11684\,
            PADOUT => \N__11683\,
            PADIN => \N__11682\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11675\,
            DIN => \N__11674\,
            DOUT => \N__11673\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11675\,
            PADOUT => \N__11674\,
            PADIN => \N__11673\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6319\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11666\,
            DIN => \N__11665\,
            DOUT => \N__11664\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11666\,
            PADOUT => \N__11665\,
            PADIN => \N__11664\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6148\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11657\,
            DIN => \N__11656\,
            DOUT => \N__11655\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11657\,
            PADOUT => \N__11656\,
            PADIN => \N__11655\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9077\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11648\,
            DIN => \N__11647\,
            DOUT => \N__11646\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11648\,
            PADOUT => \N__11647\,
            PADIN => \N__11646\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4147\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11639\,
            DIN => \N__11638\,
            DOUT => \N__11637\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11639\,
            PADOUT => \N__11638\,
            PADIN => \N__11637\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11630\,
            DIN => \N__11629\,
            DOUT => \N__11628\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11630\,
            PADOUT => \N__11629\,
            PADIN => \N__11628\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8890\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11621\,
            DIN => \N__11620\,
            DOUT => \N__11619\,
            PACKAGEPIN => \DA_wire\(0)
        );

    \DA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11621\,
            PADOUT => \N__11620\,
            PADIN => \N__11619\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4990\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11612\,
            DIN => \N__11611\,
            DOUT => \N__11610\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11612\,
            PADOUT => \N__11611\,
            PADIN => \N__11610\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7954\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11603\,
            DIN => \N__11602\,
            DOUT => \N__11601\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11603\,
            PADOUT => \N__11602\,
            PADIN => \N__11601\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11594\,
            DIN => \N__11593\,
            DOUT => \N__11592\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11594\,
            PADOUT => \N__11593\,
            PADIN => \N__11592\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11585\,
            DIN => \N__11584\,
            DOUT => \N__11583\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11585\,
            PADOUT => \N__11584\,
            PADIN => \N__11583\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11576\,
            DIN => \N__11575\,
            DOUT => \N__11574\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11576\,
            PADOUT => \N__11575\,
            PADIN => \N__11574\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11567\,
            DIN => \N__11566\,
            DOUT => \N__11565\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11567\,
            PADOUT => \N__11566\,
            PADIN => \N__11565\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7588\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11558\,
            DIN => \N__11557\,
            DOUT => \N__11556\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11558\,
            PADOUT => \N__11557\,
            PADIN => \N__11556\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11549\,
            DIN => \N__11548\,
            DOUT => \N__11547\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11549\,
            PADOUT => \N__11548\,
            PADIN => \N__11547\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9081\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11540\,
            DIN => \N__11539\,
            DOUT => \N__11538\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11540\,
            PADOUT => \N__11539\,
            PADIN => \N__11538\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11531\,
            DIN => \N__11530\,
            DOUT => \N__11529\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11531\,
            PADOUT => \N__11530\,
            PADIN => \N__11529\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11038\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11522\,
            DIN => \N__11521\,
            DOUT => \N__11520\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11522\,
            PADOUT => \N__11521\,
            PADIN => \N__11520\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9154\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11513\,
            DIN => \N__11512\,
            DOUT => \N__11511\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11513\,
            PADOUT => \N__11512\,
            PADIN => \N__11511\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6289\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11504\,
            DIN => \N__11503\,
            DOUT => \N__11502\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11504\,
            PADOUT => \N__11503\,
            PADIN => \N__11502\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4564\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11495\,
            DIN => \N__11494\,
            DOUT => \N__11493\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11495\,
            PADOUT => \N__11494\,
            PADIN => \N__11493\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11486\,
            DIN => \N__11485\,
            DOUT => \N__11484\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11486\,
            PADOUT => \N__11485\,
            PADIN => \N__11484\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11477\,
            DIN => \N__11476\,
            DOUT => \N__11475\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11477\,
            PADOUT => \N__11476\,
            PADIN => \N__11475\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7858\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11468\,
            DIN => \N__11467\,
            DOUT => \N__11466\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11468\,
            PADOUT => \N__11467\,
            PADIN => \N__11466\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4709\,
            DIN0 => OPEN,
            DOUT0 => \N__4633\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11459\,
            DIN => \N__11458\,
            DOUT => \N__11457\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11459\,
            PADOUT => \N__11458\,
            PADIN => \N__11457\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9796\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11450\,
            DIN => \N__11449\,
            DOUT => \N__11448\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11450\,
            PADOUT => \N__11449\,
            PADIN => \N__11448\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4180\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11441\,
            DIN => \N__11440\,
            DOUT => \N__11439\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11441\,
            PADOUT => \N__11440\,
            PADIN => \N__11439\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7006\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11432\,
            DIN => \N__11431\,
            DOUT => \N__11430\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11432\,
            PADOUT => \N__11431\,
            PADIN => \N__11430\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11423\,
            DIN => \N__11422\,
            DOUT => \N__11421\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11423\,
            PADOUT => \N__11422\,
            PADIN => \N__11421\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11414\,
            DIN => \N__11413\,
            DOUT => \N__11412\,
            PACKAGEPIN => \DA_wire\(2)
        );

    \DA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11414\,
            PADOUT => \N__11413\,
            PADIN => \N__11412\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11405\,
            DIN => \N__11404\,
            DOUT => \N__11403\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11405\,
            PADOUT => \N__11404\,
            PADIN => \N__11403\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11396\,
            DIN => \N__11395\,
            DOUT => \N__11394\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11396\,
            PADOUT => \N__11395\,
            PADIN => \N__11394\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11387\,
            DIN => \N__11386\,
            DOUT => \N__11385\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11387\,
            PADOUT => \N__11386\,
            PADIN => \N__11385\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7600\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11378\,
            DIN => \N__11377\,
            DOUT => \N__11376\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11378\,
            PADOUT => \N__11377\,
            PADIN => \N__11376\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8281\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11369\,
            DIN => \N__11368\,
            DOUT => \N__11367\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11369\,
            PADOUT => \N__11368\,
            PADIN => \N__11367\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11360\,
            DIN => \N__11359\,
            DOUT => \N__11358\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11360\,
            PADOUT => \N__11359\,
            PADIN => \N__11358\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11351\,
            DIN => \N__11350\,
            DOUT => \N__11349\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11351\,
            PADOUT => \N__11350\,
            PADIN => \N__11349\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4710\,
            DIN0 => OPEN,
            DOUT0 => \N__4622\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11342\,
            DIN => \N__11341\,
            DOUT => \N__11340\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11342\,
            PADOUT => \N__11341\,
            PADIN => \N__11340\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8065\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11333\,
            DIN => \N__11332\,
            DOUT => \N__11331\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11333\,
            PADOUT => \N__11332\,
            PADIN => \N__11331\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11324\,
            DIN => \N__11323\,
            DOUT => \N__11322\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11324\,
            PADOUT => \N__11323\,
            PADIN => \N__11322\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11315\,
            DIN => \N__11314\,
            DOUT => \N__11313\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11315\,
            PADOUT => \N__11314\,
            PADIN => \N__11313\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11306\,
            DIN => \N__11305\,
            DOUT => \N__11304\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11306\,
            PADOUT => \N__11305\,
            PADIN => \N__11304\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11297\,
            DIN => \N__11296\,
            DOUT => \N__11295\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11297\,
            PADOUT => \N__11296\,
            PADIN => \N__11295\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11288\,
            DIN => \N__11287\,
            DOUT => \N__11286\,
            PACKAGEPIN => \DA_wire\(1)
        );

    \DA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11288\,
            PADOUT => \N__11287\,
            PADIN => \N__11286\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7516\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11279\,
            DIN => \N__11278\,
            DOUT => \N__11277\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11279\,
            PADOUT => \N__11278\,
            PADIN => \N__11277\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11270\,
            DIN => \N__11269\,
            DOUT => \N__11268\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11270\,
            PADOUT => \N__11269\,
            PADIN => \N__11268\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11261\,
            DIN => \N__11260\,
            DOUT => \N__11259\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11261\,
            PADOUT => \N__11260\,
            PADIN => \N__11259\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11252\,
            DIN => \N__11251\,
            DOUT => \N__11250\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11252\,
            PADOUT => \N__11251\,
            PADIN => \N__11250\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6349\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11243\,
            DIN => \N__11242\,
            DOUT => \N__11241\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11243\,
            PADOUT => \N__11242\,
            PADIN => \N__11241\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8623\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11234\,
            DIN => \N__11233\,
            DOUT => \N__11232\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11234\,
            PADOUT => \N__11233\,
            PADIN => \N__11232\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4333\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11225\,
            DIN => \N__11224\,
            DOUT => \N__11223\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11225\,
            PADOUT => \N__11224\,
            PADIN => \N__11223\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11216\,
            DIN => \N__11215\,
            DOUT => \N__11214\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11216\,
            PADOUT => \N__11215\,
            PADIN => \N__11214\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11207\,
            DIN => \N__11206\,
            DOUT => \N__11205\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11207\,
            PADOUT => \N__11206\,
            PADIN => \N__11205\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7567\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11198\,
            DIN => \N__11197\,
            DOUT => \N__11196\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11198\,
            PADOUT => \N__11197\,
            PADIN => \N__11196\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11189\,
            DIN => \N__11188\,
            DOUT => \N__11187\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11189\,
            PADOUT => \N__11188\,
            PADIN => \N__11187\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11180\,
            DIN => \N__11179\,
            DOUT => \N__11178\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11180\,
            PADOUT => \N__11179\,
            PADIN => \N__11178\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6664\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11171\,
            DIN => \N__11170\,
            DOUT => \N__11169\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11171\,
            PADOUT => \N__11170\,
            PADIN => \N__11169\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11162\,
            DIN => \N__11161\,
            DOUT => \N__11160\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11162\,
            PADOUT => \N__11161\,
            PADIN => \N__11160\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9085\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11153\,
            DIN => \N__11152\,
            DOUT => \N__11151\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11153\,
            PADOUT => \N__11152\,
            PADIN => \N__11151\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2710\ : InMux
    port map (
            O => \N__11134\,
            I => \N__11129\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11133\,
            I => \N__11124\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11132\,
            I => \N__11124\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11129\,
            I => \N__11118\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11118\
        );

    \I__2705\ : InMux
    port map (
            O => \N__11123\,
            I => \N__11115\
        );

    \I__2704\ : Span4Mux_v
    port map (
            O => \N__11118\,
            I => \N__11112\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__11115\,
            I => \N__11109\
        );

    \I__2702\ : Span4Mux_v
    port map (
            O => \N__11112\,
            I => \N__11104\
        );

    \I__2701\ : Span4Mux_h
    port map (
            O => \N__11109\,
            I => \N__11104\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__11104\,
            I => \N__11100\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11096\
        );

    \I__2698\ : Span4Mux_h
    port map (
            O => \N__11100\,
            I => \N__11093\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11099\,
            I => \N__11088\
        );

    \I__2696\ : InMux
    port map (
            O => \N__11096\,
            I => \N__11088\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__11093\,
            I => \N__11083\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__11088\,
            I => \N__11083\
        );

    \I__2693\ : Span4Mux_h
    port map (
            O => \N__11083\,
            I => \N__11080\
        );

    \I__2692\ : Span4Mux_v
    port map (
            O => \N__11080\,
            I => \N__11077\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__11077\,
            I => \CASUn_c\
        );

    \I__2690\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11071\,
            I => \N__11068\
        );

    \I__2688\ : Span4Mux_v
    port map (
            O => \N__11068\,
            I => \N__11064\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11067\,
            I => \N__11061\
        );

    \I__2686\ : Sp12to4
    port map (
            O => \N__11064\,
            I => \N__11058\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11055\
        );

    \I__2684\ : Span12Mux_h
    port map (
            O => \N__11058\,
            I => \N__11051\
        );

    \I__2683\ : Sp12to4
    port map (
            O => \N__11055\,
            I => \N__11048\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11045\
        );

    \I__2681\ : Odrv12
    port map (
            O => \N__11051\,
            I => \REG_CYCLEm\
        );

    \I__2680\ : Odrv12
    port map (
            O => \N__11048\,
            I => \REG_CYCLEm\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11045\,
            I => \REG_CYCLEm\
        );

    \I__2678\ : IoInMux
    port map (
            O => \N__11038\,
            I => \N__11035\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11035\,
            I => \N__11032\
        );

    \I__2676\ : Span4Mux_s3_v
    port map (
            O => \N__11032\,
            I => \N__11029\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__11029\,
            I => \N__11026\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__11026\,
            I => \DRDENn_c\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11023\,
            I => \N__11020\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__11020\,
            I => \N__11015\
        );

    \I__2671\ : InMux
    port map (
            O => \N__11019\,
            I => \N__11012\
        );

    \I__2670\ : InMux
    port map (
            O => \N__11018\,
            I => \N__11009\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__11015\,
            I => \N__11005\
        );

    \I__2668\ : LocalMux
    port map (
            O => \N__11012\,
            I => \N__11000\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__11009\,
            I => \N__11000\
        );

    \I__2666\ : InMux
    port map (
            O => \N__11008\,
            I => \N__10997\
        );

    \I__2665\ : Sp12to4
    port map (
            O => \N__11005\,
            I => \N__10990\
        );

    \I__2664\ : Sp12to4
    port map (
            O => \N__11000\,
            I => \N__10990\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__10997\,
            I => \N__10990\
        );

    \I__2662\ : Span12Mux_v
    port map (
            O => \N__10990\,
            I => \N__10987\
        );

    \I__2661\ : Span12Mux_h
    port map (
            O => \N__10987\,
            I => \N__10984\
        );

    \I__2660\ : Odrv12
    port map (
            O => \N__10984\,
            I => \DRA_c_1\
        );

    \I__2659\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10977\
        );

    \I__2658\ : InMux
    port map (
            O => \N__10980\,
            I => \N__10974\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10971\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10968\
        );

    \I__2655\ : Span4Mux_h
    port map (
            O => \N__10971\,
            I => \N__10963\
        );

    \I__2654\ : Span4Mux_v
    port map (
            O => \N__10968\,
            I => \N__10963\
        );

    \I__2653\ : Sp12to4
    port map (
            O => \N__10963\,
            I => \N__10960\
        );

    \I__2652\ : Span12Mux_h
    port map (
            O => \N__10960\,
            I => \N__10957\
        );

    \I__2651\ : Span12Mux_v
    port map (
            O => \N__10957\,
            I => \N__10954\
        );

    \I__2650\ : Odrv12
    port map (
            O => \N__10954\,
            I => \DRA_c_0\
        );

    \I__2649\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10948\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10945\
        );

    \I__2647\ : Span4Mux_h
    port map (
            O => \N__10945\,
            I => \N__10942\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__10942\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__2645\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10934\
        );

    \I__2644\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10931\
        );

    \I__2643\ : InMux
    port map (
            O => \N__10937\,
            I => \N__10928\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10920\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10920\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10920\
        );

    \I__2639\ : InMux
    port map (
            O => \N__10927\,
            I => \N__10917\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__10920\,
            I => \N__10914\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10911\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__10914\,
            I => \N__10908\
        );

    \I__2635\ : Sp12to4
    port map (
            O => \N__10911\,
            I => \N__10905\
        );

    \I__2634\ : Sp12to4
    port map (
            O => \N__10908\,
            I => \N__10900\
        );

    \I__2633\ : Span12Mux_v
    port map (
            O => \N__10905\,
            I => \N__10900\
        );

    \I__2632\ : Span12Mux_h
    port map (
            O => \N__10900\,
            I => \N__10897\
        );

    \I__2631\ : Odrv12
    port map (
            O => \N__10897\,
            I => \DRA_c_4\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10894\,
            I => \N__10887\
        );

    \I__2629\ : InMux
    port map (
            O => \N__10893\,
            I => \N__10887\
        );

    \I__2628\ : InMux
    port map (
            O => \N__10892\,
            I => \N__10883\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__10887\,
            I => \N__10880\
        );

    \I__2626\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10877\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10870\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10870\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__10877\,
            I => \N__10870\
        );

    \I__2622\ : Span4Mux_h
    port map (
            O => \N__10870\,
            I => \N__10867\
        );

    \I__2621\ : Sp12to4
    port map (
            O => \N__10867\,
            I => \N__10864\
        );

    \I__2620\ : Span12Mux_v
    port map (
            O => \N__10864\,
            I => \N__10861\
        );

    \I__2619\ : Odrv12
    port map (
            O => \N__10861\,
            I => \DRA_c_3\
        );

    \I__2618\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10855\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__10855\,
            I => \N__10852\
        );

    \I__2616\ : Odrv12
    port map (
            O => \N__10852\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__10849\,
            I => \N__10846\
        );

    \I__2614\ : InMux
    port map (
            O => \N__10846\,
            I => \N__10843\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__10843\,
            I => \N__10840\
        );

    \I__2612\ : Span4Mux_v
    port map (
            O => \N__10840\,
            I => \N__10837\
        );

    \I__2611\ : Odrv4
    port map (
            O => \N__10837\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__2610\ : InMux
    port map (
            O => \N__10834\,
            I => \N__10828\
        );

    \I__2609\ : InMux
    port map (
            O => \N__10833\,
            I => \N__10825\
        );

    \I__2608\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10820\
        );

    \I__2607\ : InMux
    port map (
            O => \N__10831\,
            I => \N__10820\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__10828\,
            I => \N__10817\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__10825\,
            I => \N__10812\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10812\
        );

    \I__2603\ : Span4Mux_v
    port map (
            O => \N__10817\,
            I => \N__10809\
        );

    \I__2602\ : Span4Mux_v
    port map (
            O => \N__10812\,
            I => \N__10806\
        );

    \I__2601\ : Sp12to4
    port map (
            O => \N__10809\,
            I => \N__10801\
        );

    \I__2600\ : Sp12to4
    port map (
            O => \N__10806\,
            I => \N__10801\
        );

    \I__2599\ : Span12Mux_h
    port map (
            O => \N__10801\,
            I => \N__10798\
        );

    \I__2598\ : Odrv12
    port map (
            O => \N__10798\,
            I => \DRA_c_8\
        );

    \I__2597\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10792\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10789\
        );

    \I__2595\ : Span4Mux_h
    port map (
            O => \N__10789\,
            I => \N__10786\
        );

    \I__2594\ : Odrv4
    port map (
            O => \N__10786\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10776\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10782\,
            I => \N__10776\
        );

    \I__2591\ : InMux
    port map (
            O => \N__10781\,
            I => \N__10773\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10776\,
            I => \N__10767\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__2588\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10764\
        );

    \I__2587\ : Span4Mux_v
    port map (
            O => \N__10767\,
            I => \N__10761\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__2585\ : Span4Mux_h
    port map (
            O => \N__10761\,
            I => \N__10753\
        );

    \I__2584\ : Span4Mux_v
    port map (
            O => \N__10758\,
            I => \N__10753\
        );

    \I__2583\ : Sp12to4
    port map (
            O => \N__10753\,
            I => \N__10750\
        );

    \I__2582\ : Odrv12
    port map (
            O => \N__10750\,
            I => \DRA_c_6\
        );

    \I__2581\ : InMux
    port map (
            O => \N__10747\,
            I => \N__10741\
        );

    \I__2580\ : InMux
    port map (
            O => \N__10746\,
            I => \N__10738\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10735\
        );

    \I__2578\ : InMux
    port map (
            O => \N__10744\,
            I => \N__10732\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__10741\,
            I => \N__10725\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__10738\,
            I => \N__10725\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__10735\,
            I => \N__10725\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10722\
        );

    \I__2573\ : Span12Mux_h
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__2572\ : Span12Mux_h
    port map (
            O => \N__10722\,
            I => \N__10716\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__10719\,
            I => \DRA_c_7\
        );

    \I__2570\ : Odrv12
    port map (
            O => \N__10716\,
            I => \DRA_c_7\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10711\,
            I => \N__10708\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__10708\,
            I => \N__10705\
        );

    \I__2567\ : Span4Mux_h
    port map (
            O => \N__10705\,
            I => \N__10702\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__10702\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__2565\ : CascadeMux
    port map (
            O => \N__10699\,
            I => \N__10694\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10690\
        );

    \I__2563\ : CascadeMux
    port map (
            O => \N__10697\,
            I => \N__10682\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10675\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10693\,
            I => \N__10670\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__10690\,
            I => \N__10662\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10659\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10688\,
            I => \N__10654\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10687\,
            I => \N__10654\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10645\
        );

    \I__2555\ : InMux
    port map (
            O => \N__10685\,
            I => \N__10645\
        );

    \I__2554\ : InMux
    port map (
            O => \N__10682\,
            I => \N__10645\
        );

    \I__2553\ : InMux
    port map (
            O => \N__10681\,
            I => \N__10645\
        );

    \I__2552\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10642\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10637\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10637\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10634\
        );

    \I__2548\ : InMux
    port map (
            O => \N__10674\,
            I => \N__10629\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10629\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__10670\,
            I => \N__10626\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10623\
        );

    \I__2544\ : InMux
    port map (
            O => \N__10668\,
            I => \N__10620\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10667\,
            I => \N__10613\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10613\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10613\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__10662\,
            I => \N__10610\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__10659\,
            I => \N__10599\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10654\,
            I => \N__10599\
        );

    \I__2537\ : LocalMux
    port map (
            O => \N__10645\,
            I => \N__10599\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10599\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__10637\,
            I => \N__10599\
        );

    \I__2534\ : Span4Mux_v
    port map (
            O => \N__10634\,
            I => \N__10593\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10629\,
            I => \N__10593\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__10626\,
            I => \N__10586\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10623\,
            I => \N__10586\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10620\,
            I => \N__10586\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10613\,
            I => \N__10583\
        );

    \I__2528\ : Span4Mux_h
    port map (
            O => \N__10610\,
            I => \N__10578\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__10599\,
            I => \N__10578\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10598\,
            I => \N__10575\
        );

    \I__2525\ : Span4Mux_h
    port map (
            O => \N__10593\,
            I => \N__10570\
        );

    \I__2524\ : Span4Mux_v
    port map (
            O => \N__10586\,
            I => \N__10570\
        );

    \I__2523\ : Sp12to4
    port map (
            O => \N__10583\,
            I => \N__10567\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__10578\,
            I => \N__10560\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10575\,
            I => \N__10560\
        );

    \I__2520\ : Sp12to4
    port map (
            O => \N__10570\,
            I => \N__10560\
        );

    \I__2519\ : Span12Mux_v
    port map (
            O => \N__10567\,
            I => \N__10557\
        );

    \I__2518\ : Span12Mux_h
    port map (
            O => \N__10560\,
            I => \N__10554\
        );

    \I__2517\ : Span12Mux_h
    port map (
            O => \N__10557\,
            I => \N__10549\
        );

    \I__2516\ : Span12Mux_v
    port map (
            O => \N__10554\,
            I => \N__10549\
        );

    \I__2515\ : Odrv12
    port map (
            O => \N__10549\,
            I => \AGNUS_REV_c\
        );

    \I__2514\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10541\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10538\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10534\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__10541\,
            I => \N__10529\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10538\,
            I => \N__10529\
        );

    \I__2509\ : InMux
    port map (
            O => \N__10537\,
            I => \N__10526\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10523\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__10529\,
            I => \N__10518\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__10526\,
            I => \N__10518\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__10523\,
            I => \N__10513\
        );

    \I__2504\ : Span4Mux_h
    port map (
            O => \N__10518\,
            I => \N__10513\
        );

    \I__2503\ : Sp12to4
    port map (
            O => \N__10513\,
            I => \N__10510\
        );

    \I__2502\ : Span12Mux_v
    port map (
            O => \N__10510\,
            I => \N__10507\
        );

    \I__2501\ : Odrv12
    port map (
            O => \N__10507\,
            I => \DRA_c_9\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10501\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10501\,
            I => \N__10498\
        );

    \I__2498\ : Span12Mux_h
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__2497\ : Odrv12
    port map (
            O => \N__10495\,
            I => \RAS0n_c\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10492\,
            I => \N__10489\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__10489\,
            I => \N__10486\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__10486\,
            I => \N__10483\
        );

    \I__2493\ : Span4Mux_h
    port map (
            O => \N__10483\,
            I => \N__10480\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__10480\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2491\ : ClkMux
    port map (
            O => \N__10477\,
            I => \N__10462\
        );

    \I__2490\ : ClkMux
    port map (
            O => \N__10476\,
            I => \N__10462\
        );

    \I__2489\ : ClkMux
    port map (
            O => \N__10475\,
            I => \N__10462\
        );

    \I__2488\ : ClkMux
    port map (
            O => \N__10474\,
            I => \N__10462\
        );

    \I__2487\ : ClkMux
    port map (
            O => \N__10473\,
            I => \N__10462\
        );

    \I__2486\ : GlobalMux
    port map (
            O => \N__10462\,
            I => \N__10459\
        );

    \I__2485\ : gio2CtrlBuf
    port map (
            O => \N__10459\,
            I => \C3_c_g\
        );

    \I__2484\ : CEMux
    port map (
            O => \N__10456\,
            I => \N__10423\
        );

    \I__2483\ : CEMux
    port map (
            O => \N__10455\,
            I => \N__10423\
        );

    \I__2482\ : CEMux
    port map (
            O => \N__10454\,
            I => \N__10423\
        );

    \I__2481\ : CEMux
    port map (
            O => \N__10453\,
            I => \N__10423\
        );

    \I__2480\ : CEMux
    port map (
            O => \N__10452\,
            I => \N__10423\
        );

    \I__2479\ : CEMux
    port map (
            O => \N__10451\,
            I => \N__10423\
        );

    \I__2478\ : CEMux
    port map (
            O => \N__10450\,
            I => \N__10423\
        );

    \I__2477\ : CEMux
    port map (
            O => \N__10449\,
            I => \N__10423\
        );

    \I__2476\ : CEMux
    port map (
            O => \N__10448\,
            I => \N__10423\
        );

    \I__2475\ : CEMux
    port map (
            O => \N__10447\,
            I => \N__10423\
        );

    \I__2474\ : CEMux
    port map (
            O => \N__10446\,
            I => \N__10423\
        );

    \I__2473\ : GlobalMux
    port map (
            O => \N__10423\,
            I => \N__10420\
        );

    \I__2472\ : gio2CtrlBuf
    port map (
            O => \N__10420\,
            I => \DBRn_c_i_0_g\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10410\
        );

    \I__2470\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10407\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10402\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10414\,
            I => \N__10402\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10399\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10410\,
            I => \N__10396\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__10407\,
            I => \N__10380\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10402\,
            I => \N__10377\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10399\,
            I => \N__10356\
        );

    \I__2462\ : Glb2LocalMux
    port map (
            O => \N__10396\,
            I => \N__10276\
        );

    \I__2461\ : SRMux
    port map (
            O => \N__10395\,
            I => \N__10276\
        );

    \I__2460\ : SRMux
    port map (
            O => \N__10394\,
            I => \N__10276\
        );

    \I__2459\ : SRMux
    port map (
            O => \N__10393\,
            I => \N__10276\
        );

    \I__2458\ : SRMux
    port map (
            O => \N__10392\,
            I => \N__10276\
        );

    \I__2457\ : SRMux
    port map (
            O => \N__10391\,
            I => \N__10276\
        );

    \I__2456\ : SRMux
    port map (
            O => \N__10390\,
            I => \N__10276\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__10389\,
            I => \N__10276\
        );

    \I__2454\ : SRMux
    port map (
            O => \N__10388\,
            I => \N__10276\
        );

    \I__2453\ : SRMux
    port map (
            O => \N__10387\,
            I => \N__10276\
        );

    \I__2452\ : SRMux
    port map (
            O => \N__10386\,
            I => \N__10276\
        );

    \I__2451\ : SRMux
    port map (
            O => \N__10385\,
            I => \N__10276\
        );

    \I__2450\ : SRMux
    port map (
            O => \N__10384\,
            I => \N__10276\
        );

    \I__2449\ : SRMux
    port map (
            O => \N__10383\,
            I => \N__10276\
        );

    \I__2448\ : Glb2LocalMux
    port map (
            O => \N__10380\,
            I => \N__10276\
        );

    \I__2447\ : Glb2LocalMux
    port map (
            O => \N__10377\,
            I => \N__10276\
        );

    \I__2446\ : SRMux
    port map (
            O => \N__10376\,
            I => \N__10276\
        );

    \I__2445\ : SRMux
    port map (
            O => \N__10375\,
            I => \N__10276\
        );

    \I__2444\ : SRMux
    port map (
            O => \N__10374\,
            I => \N__10276\
        );

    \I__2443\ : SRMux
    port map (
            O => \N__10373\,
            I => \N__10276\
        );

    \I__2442\ : SRMux
    port map (
            O => \N__10372\,
            I => \N__10276\
        );

    \I__2441\ : SRMux
    port map (
            O => \N__10371\,
            I => \N__10276\
        );

    \I__2440\ : SRMux
    port map (
            O => \N__10370\,
            I => \N__10276\
        );

    \I__2439\ : SRMux
    port map (
            O => \N__10369\,
            I => \N__10276\
        );

    \I__2438\ : SRMux
    port map (
            O => \N__10368\,
            I => \N__10276\
        );

    \I__2437\ : SRMux
    port map (
            O => \N__10367\,
            I => \N__10276\
        );

    \I__2436\ : SRMux
    port map (
            O => \N__10366\,
            I => \N__10276\
        );

    \I__2435\ : SRMux
    port map (
            O => \N__10365\,
            I => \N__10276\
        );

    \I__2434\ : SRMux
    port map (
            O => \N__10364\,
            I => \N__10276\
        );

    \I__2433\ : SRMux
    port map (
            O => \N__10363\,
            I => \N__10276\
        );

    \I__2432\ : SRMux
    port map (
            O => \N__10362\,
            I => \N__10276\
        );

    \I__2431\ : SRMux
    port map (
            O => \N__10361\,
            I => \N__10276\
        );

    \I__2430\ : SRMux
    port map (
            O => \N__10360\,
            I => \N__10276\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__10359\,
            I => \N__10276\
        );

    \I__2428\ : Glb2LocalMux
    port map (
            O => \N__10356\,
            I => \N__10276\
        );

    \I__2427\ : SRMux
    port map (
            O => \N__10355\,
            I => \N__10276\
        );

    \I__2426\ : SRMux
    port map (
            O => \N__10354\,
            I => \N__10276\
        );

    \I__2425\ : SRMux
    port map (
            O => \N__10353\,
            I => \N__10276\
        );

    \I__2424\ : GlobalMux
    port map (
            O => \N__10276\,
            I => \N__10273\
        );

    \I__2423\ : gio2CtrlBuf
    port map (
            O => \N__10273\,
            I => \RESETn_c_i_g\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10270\,
            I => \N__10266\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10266\,
            I => \N__10257\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10263\,
            I => \N__10254\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10262\,
            I => \N__10251\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10261\,
            I => \N__10248\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10260\,
            I => \N__10245\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__10257\,
            I => \N__10242\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__10254\,
            I => \N__10237\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__10251\,
            I => \N__10237\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10248\,
            I => \N__10234\
        );

    \I__2411\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10231\
        );

    \I__2410\ : Sp12to4
    port map (
            O => \N__10242\,
            I => \N__10228\
        );

    \I__2409\ : Span4Mux_v
    port map (
            O => \N__10237\,
            I => \N__10225\
        );

    \I__2408\ : Span4Mux_v
    port map (
            O => \N__10234\,
            I => \N__10222\
        );

    \I__2407\ : Span12Mux_v
    port map (
            O => \N__10231\,
            I => \N__10219\
        );

    \I__2406\ : Span12Mux_h
    port map (
            O => \N__10228\,
            I => \N__10212\
        );

    \I__2405\ : Sp12to4
    port map (
            O => \N__10225\,
            I => \N__10212\
        );

    \I__2404\ : Sp12to4
    port map (
            O => \N__10222\,
            I => \N__10212\
        );

    \I__2403\ : Span12Mux_h
    port map (
            O => \N__10219\,
            I => \N__10209\
        );

    \I__2402\ : Span12Mux_h
    port map (
            O => \N__10212\,
            I => \N__10206\
        );

    \I__2401\ : Odrv12
    port map (
            O => \N__10209\,
            I => \RnW_c\
        );

    \I__2400\ : Odrv12
    port map (
            O => \N__10206\,
            I => \RnW_c\
        );

    \I__2399\ : InMux
    port map (
            O => \N__10201\,
            I => \N__10197\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__10200\,
            I => \N__10192\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10197\,
            I => \N__10189\
        );

    \I__2396\ : InMux
    port map (
            O => \N__10196\,
            I => \N__10186\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__10195\,
            I => \N__10182\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10192\,
            I => \N__10179\
        );

    \I__2393\ : Span12Mux_s6_h
    port map (
            O => \N__10189\,
            I => \N__10174\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10186\,
            I => \N__10174\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10168\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10168\
        );

    \I__2389\ : LocalMux
    port map (
            O => \N__10179\,
            I => \N__10164\
        );

    \I__2388\ : Span12Mux_h
    port map (
            O => \N__10174\,
            I => \N__10159\
        );

    \I__2387\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10156\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10168\,
            I => \N__10153\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10150\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__10164\,
            I => \N__10147\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10163\,
            I => \N__10142\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10162\,
            I => \N__10142\
        );

    \I__2381\ : Odrv12
    port map (
            O => \N__10159\,
            I => \WRITE_CYCLEm\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10156\,
            I => \WRITE_CYCLEm\
        );

    \I__2379\ : Odrv4
    port map (
            O => \N__10153\,
            I => \WRITE_CYCLEm\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10150\,
            I => \WRITE_CYCLEm\
        );

    \I__2377\ : Odrv4
    port map (
            O => \N__10147\,
            I => \WRITE_CYCLEm\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__10142\,
            I => \WRITE_CYCLEm\
        );

    \I__2375\ : IoInMux
    port map (
            O => \N__10129\,
            I => \N__10126\
        );

    \I__2374\ : LocalMux
    port map (
            O => \N__10126\,
            I => \N__10123\
        );

    \I__2373\ : Span4Mux_s3_h
    port map (
            O => \N__10123\,
            I => \N__10120\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__10120\,
            I => \N__10117\
        );

    \I__2371\ : Odrv4
    port map (
            O => \N__10117\,
            I => \N_405\
        );

    \I__2370\ : InMux
    port map (
            O => \N__10114\,
            I => \N__10110\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10113\,
            I => \N__10107\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__10110\,
            I => \N__10102\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__10107\,
            I => \N__10102\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__10102\,
            I => \N__10098\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10101\,
            I => \N__10095\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__10098\,
            I => \N__10090\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10095\,
            I => \N__10090\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__10090\,
            I => \N__10086\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10089\,
            I => \N__10083\
        );

    \I__2360\ : Sp12to4
    port map (
            O => \N__10086\,
            I => \N__10078\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10083\,
            I => \N__10075\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10082\,
            I => \N__10070\
        );

    \I__2357\ : InMux
    port map (
            O => \N__10081\,
            I => \N__10070\
        );

    \I__2356\ : Span12Mux_s2_v
    port map (
            O => \N__10078\,
            I => \N__10067\
        );

    \I__2355\ : Span12Mux_h
    port map (
            O => \N__10075\,
            I => \N__10062\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10070\,
            I => \N__10062\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__10067\,
            I => \N__10057\
        );

    \I__2352\ : Span12Mux_v
    port map (
            O => \N__10062\,
            I => \N__10057\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__10057\,
            I => \CASLn_c\
        );

    \I__2350\ : InMux
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__10051\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10048\,
            I => \N__10045\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__10045\,
            I => \N__10042\
        );

    \I__2346\ : Span4Mux_h
    port map (
            O => \N__10042\,
            I => \N__10039\
        );

    \I__2345\ : Odrv4
    port map (
            O => \N__10039\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10033\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10033\,
            I => \N__10030\
        );

    \I__2342\ : Odrv4
    port map (
            O => \N__10030\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2341\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10024\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__2339\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10015\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10022\,
            I => \N__10012\
        );

    \I__2337\ : InMux
    port map (
            O => \N__10021\,
            I => \N__10009\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__10018\,
            I => \N__10004\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__10004\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__10012\,
            I => \N__9999\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__9999\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__10004\,
            I => \N__9996\
        );

    \I__2331\ : Span12Mux_v
    port map (
            O => \N__9999\,
            I => \N__9991\
        );

    \I__2330\ : Sp12to4
    port map (
            O => \N__9996\,
            I => \N__9991\
        );

    \I__2329\ : Span12Mux_h
    port map (
            O => \N__9991\,
            I => \N__9988\
        );

    \I__2328\ : Odrv12
    port map (
            O => \N__9988\,
            I => \DRA_c_5\
        );

    \I__2327\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9982\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__9982\,
            I => \N__9979\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__9979\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9973\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__9973\,
            I => \N__9970\
        );

    \I__2322\ : Odrv4
    port map (
            O => \N__9970\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__2321\ : InMux
    port map (
            O => \N__9967\,
            I => \N__9964\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9964\,
            I => \N__9961\
        );

    \I__2319\ : Odrv12
    port map (
            O => \N__9961\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9958\,
            I => \N__9955\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9955\,
            I => \N__9952\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__9952\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9941\
        );

    \I__2314\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9941\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9938\
        );

    \I__2312\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9935\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__9941\,
            I => \N__9930\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__9938\,
            I => \N__9930\
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__9935\,
            I => \N__9925\
        );

    \I__2308\ : Sp12to4
    port map (
            O => \N__9930\,
            I => \N__9925\
        );

    \I__2307\ : Span12Mux_v
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__2306\ : Span12Mux_h
    port map (
            O => \N__9922\,
            I => \N__9919\
        );

    \I__2305\ : Odrv12
    port map (
            O => \N__9919\,
            I => \DRA_c_2\
        );

    \I__2304\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9913\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__2301\ : Odrv4
    port map (
            O => \N__9907\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__9904\,
            I => \N__9901\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9898\,
            I => \N__9895\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__9895\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2296\ : InMux
    port map (
            O => \N__9892\,
            I => \N__9888\
        );

    \I__2295\ : InMux
    port map (
            O => \N__9891\,
            I => \N__9885\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9882\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9885\,
            I => \N__9879\
        );

    \I__2292\ : Span4Mux_v
    port map (
            O => \N__9882\,
            I => \N__9873\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__9879\,
            I => \N__9873\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9868\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__9873\,
            I => \N__9865\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9862\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9871\,
            I => \N__9859\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9868\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2285\ : Odrv4
    port map (
            O => \N__9865\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__9862\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9859\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__2282\ : IoInMux
    port map (
            O => \N__9850\,
            I => \N__9847\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__9847\,
            I => \N__9844\
        );

    \I__2280\ : Span12Mux_s8_v
    port map (
            O => \N__9844\,
            I => \N__9841\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__9841\,
            I => \CRCSn_c\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9835\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__9835\,
            I => \N__9831\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9828\
        );

    \I__2275\ : Span4Mux_h
    port map (
            O => \N__9831\,
            I => \N__9821\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__9828\,
            I => \N__9821\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__9827\,
            I => \N__9817\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9826\,
            I => \N__9814\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__9821\,
            I => \N__9811\
        );

    \I__2270\ : InMux
    port map (
            O => \N__9820\,
            I => \N__9808\
        );

    \I__2269\ : InMux
    port map (
            O => \N__9817\,
            I => \N__9805\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__9814\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__9811\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__9808\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9805\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__2264\ : IoInMux
    port map (
            O => \N__9796\,
            I => \N__9793\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9790\
        );

    \I__2262\ : IoSpan4Mux
    port map (
            O => \N__9790\,
            I => \N__9787\
        );

    \I__2261\ : IoSpan4Mux
    port map (
            O => \N__9787\,
            I => \N__9784\
        );

    \I__2260\ : IoSpan4Mux
    port map (
            O => \N__9784\,
            I => \N__9781\
        );

    \I__2259\ : Span4Mux_s2_h
    port map (
            O => \N__9781\,
            I => \N__9778\
        );

    \I__2258\ : Sp12to4
    port map (
            O => \N__9778\,
            I => \N__9775\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__9775\,
            I => \WEn_c\
        );

    \I__2256\ : InMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__9769\,
            I => \N__9766\
        );

    \I__2254\ : Span4Mux_h
    port map (
            O => \N__9766\,
            I => \N__9763\
        );

    \I__2253\ : Odrv4
    port map (
            O => \N__9763\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2252\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9757\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9751\
        );

    \I__2250\ : InMux
    port map (
            O => \N__9756\,
            I => \N__9743\
        );

    \I__2249\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9740\
        );

    \I__2248\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9737\
        );

    \I__2247\ : Span4Mux_h
    port map (
            O => \N__9751\,
            I => \N__9734\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9729\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9729\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9724\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9747\,
            I => \N__9724\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9746\,
            I => \N__9721\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9743\,
            I => \N__9718\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9713\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9713\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__9734\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__9729\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9724\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9721\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__9718\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__9713\,
            I => \U712_CHIP_RAM.N_501\
        );

    \I__2232\ : InMux
    port map (
            O => \N__9700\,
            I => \N__9697\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9697\,
            I => \N__9683\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9676\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9695\,
            I => \N__9676\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9694\,
            I => \N__9676\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9693\,
            I => \N__9673\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9692\,
            I => \N__9668\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9668\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9663\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9663\
        );

    \I__2222\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9658\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9687\,
            I => \N__9658\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9655\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__9683\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9676\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__9673\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9668\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9663\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9658\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__9655\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__9640\,
            I => \N__9635\
        );

    \I__2211\ : CascadeMux
    port map (
            O => \N__9639\,
            I => \N__9631\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9626\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9626\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \N__9623\
        );

    \I__2207\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9620\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9626\,
            I => \N__9614\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9611\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__9620\,
            I => \N__9607\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9603\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9600\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__9617\,
            I => \N__9596\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__9614\,
            I => \N__9591\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__9611\,
            I => \N__9591\
        );

    \I__2198\ : InMux
    port map (
            O => \N__9610\,
            I => \N__9588\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__9607\,
            I => \N__9585\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9582\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9579\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9576\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9599\,
            I => \N__9573\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9596\,
            I => \N__9570\
        );

    \I__2191\ : Span4Mux_v
    port map (
            O => \N__9591\,
            I => \N__9567\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9588\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2189\ : Odrv4
    port map (
            O => \N__9585\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2188\ : LocalMux
    port map (
            O => \N__9582\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2187\ : Odrv4
    port map (
            O => \N__9579\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2186\ : Odrv4
    port map (
            O => \N__9576\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__9573\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__9570\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__9567\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__9550\,
            I => \N__9546\
        );

    \I__2181\ : InMux
    port map (
            O => \N__9549\,
            I => \N__9542\
        );

    \I__2180\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9539\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9545\,
            I => \N__9531\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9542\,
            I => \N__9524\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__9539\,
            I => \N__9521\
        );

    \I__2176\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9516\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9516\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9513\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9508\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9534\,
            I => \N__9508\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9531\,
            I => \N__9505\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9530\,
            I => \N__9502\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9499\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9494\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9494\
        );

    \I__2166\ : Odrv4
    port map (
            O => \N__9524\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2165\ : Odrv4
    port map (
            O => \N__9521\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9516\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__9513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__9508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__9505\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__9502\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9499\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9494\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__9475\,
            I => \N__9467\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9474\,
            I => \N__9464\
        );

    \I__2155\ : InMux
    port map (
            O => \N__9473\,
            I => \N__9457\
        );

    \I__2154\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9457\
        );

    \I__2153\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9457\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9454\
        );

    \I__2151\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9451\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__9464\,
            I => \N__9447\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9457\,
            I => \N__9444\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9454\,
            I => \N__9441\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__9451\,
            I => \N__9438\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9435\
        );

    \I__2145\ : Span4Mux_v
    port map (
            O => \N__9447\,
            I => \N__9432\
        );

    \I__2144\ : Span4Mux_v
    port map (
            O => \N__9444\,
            I => \N__9427\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__9441\,
            I => \N__9427\
        );

    \I__2142\ : Span12Mux_v
    port map (
            O => \N__9438\,
            I => \N__9422\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9435\,
            I => \N__9422\
        );

    \I__2140\ : Odrv4
    port map (
            O => \N__9432\,
            I => \DMA_CYCLEm\
        );

    \I__2139\ : Odrv4
    port map (
            O => \N__9427\,
            I => \DMA_CYCLEm\
        );

    \I__2138\ : Odrv12
    port map (
            O => \N__9422\,
            I => \DMA_CYCLEm\
        );

    \I__2137\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9412\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9412\,
            I => \N__9375\
        );

    \I__2135\ : ClkMux
    port map (
            O => \N__9411\,
            I => \N__9289\
        );

    \I__2134\ : ClkMux
    port map (
            O => \N__9410\,
            I => \N__9289\
        );

    \I__2133\ : ClkMux
    port map (
            O => \N__9409\,
            I => \N__9289\
        );

    \I__2132\ : ClkMux
    port map (
            O => \N__9408\,
            I => \N__9289\
        );

    \I__2131\ : ClkMux
    port map (
            O => \N__9407\,
            I => \N__9289\
        );

    \I__2130\ : ClkMux
    port map (
            O => \N__9406\,
            I => \N__9289\
        );

    \I__2129\ : ClkMux
    port map (
            O => \N__9405\,
            I => \N__9289\
        );

    \I__2128\ : ClkMux
    port map (
            O => \N__9404\,
            I => \N__9289\
        );

    \I__2127\ : ClkMux
    port map (
            O => \N__9403\,
            I => \N__9289\
        );

    \I__2126\ : ClkMux
    port map (
            O => \N__9402\,
            I => \N__9289\
        );

    \I__2125\ : ClkMux
    port map (
            O => \N__9401\,
            I => \N__9289\
        );

    \I__2124\ : ClkMux
    port map (
            O => \N__9400\,
            I => \N__9289\
        );

    \I__2123\ : ClkMux
    port map (
            O => \N__9399\,
            I => \N__9289\
        );

    \I__2122\ : ClkMux
    port map (
            O => \N__9398\,
            I => \N__9289\
        );

    \I__2121\ : ClkMux
    port map (
            O => \N__9397\,
            I => \N__9289\
        );

    \I__2120\ : ClkMux
    port map (
            O => \N__9396\,
            I => \N__9289\
        );

    \I__2119\ : ClkMux
    port map (
            O => \N__9395\,
            I => \N__9289\
        );

    \I__2118\ : ClkMux
    port map (
            O => \N__9394\,
            I => \N__9289\
        );

    \I__2117\ : ClkMux
    port map (
            O => \N__9393\,
            I => \N__9289\
        );

    \I__2116\ : ClkMux
    port map (
            O => \N__9392\,
            I => \N__9289\
        );

    \I__2115\ : ClkMux
    port map (
            O => \N__9391\,
            I => \N__9289\
        );

    \I__2114\ : ClkMux
    port map (
            O => \N__9390\,
            I => \N__9289\
        );

    \I__2113\ : ClkMux
    port map (
            O => \N__9389\,
            I => \N__9289\
        );

    \I__2112\ : ClkMux
    port map (
            O => \N__9388\,
            I => \N__9289\
        );

    \I__2111\ : ClkMux
    port map (
            O => \N__9387\,
            I => \N__9289\
        );

    \I__2110\ : ClkMux
    port map (
            O => \N__9386\,
            I => \N__9289\
        );

    \I__2109\ : ClkMux
    port map (
            O => \N__9385\,
            I => \N__9289\
        );

    \I__2108\ : ClkMux
    port map (
            O => \N__9384\,
            I => \N__9289\
        );

    \I__2107\ : ClkMux
    port map (
            O => \N__9383\,
            I => \N__9289\
        );

    \I__2106\ : ClkMux
    port map (
            O => \N__9382\,
            I => \N__9289\
        );

    \I__2105\ : ClkMux
    port map (
            O => \N__9381\,
            I => \N__9289\
        );

    \I__2104\ : ClkMux
    port map (
            O => \N__9380\,
            I => \N__9289\
        );

    \I__2103\ : ClkMux
    port map (
            O => \N__9379\,
            I => \N__9289\
        );

    \I__2102\ : ClkMux
    port map (
            O => \N__9378\,
            I => \N__9289\
        );

    \I__2101\ : Glb2LocalMux
    port map (
            O => \N__9375\,
            I => \N__9289\
        );

    \I__2100\ : ClkMux
    port map (
            O => \N__9374\,
            I => \N__9289\
        );

    \I__2099\ : ClkMux
    port map (
            O => \N__9373\,
            I => \N__9289\
        );

    \I__2098\ : ClkMux
    port map (
            O => \N__9372\,
            I => \N__9289\
        );

    \I__2097\ : ClkMux
    port map (
            O => \N__9371\,
            I => \N__9289\
        );

    \I__2096\ : ClkMux
    port map (
            O => \N__9370\,
            I => \N__9289\
        );

    \I__2095\ : GlobalMux
    port map (
            O => \N__9289\,
            I => \CLK80_PLL\
        );

    \I__2094\ : CEMux
    port map (
            O => \N__9286\,
            I => \N__9283\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__2092\ : Span4Mux_h
    port map (
            O => \N__9280\,
            I => \N__9277\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__9277\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9271\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9271\,
            I => \N__9268\
        );

    \I__2088\ : Span4Mux_v
    port map (
            O => \N__9268\,
            I => \N__9264\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9261\
        );

    \I__2086\ : Sp12to4
    port map (
            O => \N__9264\,
            I => \N__9256\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9261\,
            I => \N__9256\
        );

    \I__2084\ : Odrv12
    port map (
            O => \N__9256\,
            I => \DBRn_c_i\
        );

    \I__2083\ : InMux
    port map (
            O => \N__9253\,
            I => \N__9250\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9250\,
            I => \N__9246\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9249\,
            I => \N__9243\
        );

    \I__2080\ : Span4Mux_h
    port map (
            O => \N__9246\,
            I => \N__9240\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__9243\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9240\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9232\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9229\,
            I => \N__9223\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9228\,
            I => \N__9223\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__2072\ : Odrv4
    port map (
            O => \N__9220\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9214\,
            I => \N__9211\
        );

    \I__2069\ : Span4Mux_h
    port map (
            O => \N__9211\,
            I => \N__9208\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__9208\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2067\ : IoInMux
    port map (
            O => \N__9205\,
            I => \N__9202\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__2065\ : IoSpan4Mux
    port map (
            O => \N__9199\,
            I => \N__9196\
        );

    \I__2064\ : IoSpan4Mux
    port map (
            O => \N__9196\,
            I => \N__9192\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9189\
        );

    \I__2062\ : Sp12to4
    port map (
            O => \N__9192\,
            I => \N__9183\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9189\,
            I => \N__9180\
        );

    \I__2060\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9173\
        );

    \I__2059\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9173\
        );

    \I__2058\ : InMux
    port map (
            O => \N__9186\,
            I => \N__9173\
        );

    \I__2057\ : Span12Mux_s7_v
    port map (
            O => \N__9183\,
            I => \N__9165\
        );

    \I__2056\ : Sp12to4
    port map (
            O => \N__9180\,
            I => \N__9165\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__9173\,
            I => \N__9165\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9162\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__9165\,
            I => \DBENn_c\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9162\,
            I => \DBENn_c\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \U712_BYTE_ENABLE.N_453_cascade_\
        );

    \I__2050\ : IoInMux
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__2048\ : Span4Mux_s3_v
    port map (
            O => \N__9148\,
            I => \N__9145\
        );

    \I__2047\ : Span4Mux_h
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__2046\ : Sp12to4
    port map (
            O => \N__9142\,
            I => \N__9139\
        );

    \I__2045\ : Span12Mux_s10_v
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__9136\,
            I => \N_202_i\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9133\,
            I => \N__9128\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9132\,
            I => \N__9125\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__9131\,
            I => \N__9121\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9128\,
            I => \N__9118\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9125\,
            I => \N__9115\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9112\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9109\
        );

    \I__2036\ : Span4Mux_v
    port map (
            O => \N__9118\,
            I => \N__9106\
        );

    \I__2035\ : Span4Mux_h
    port map (
            O => \N__9115\,
            I => \N__9103\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9112\,
            I => \N__9098\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9109\,
            I => \N__9098\
        );

    \I__2032\ : Sp12to4
    port map (
            O => \N__9106\,
            I => \N__9091\
        );

    \I__2031\ : Sp12to4
    port map (
            O => \N__9103\,
            I => \N__9091\
        );

    \I__2030\ : Span12Mux_h
    port map (
            O => \N__9098\,
            I => \N__9091\
        );

    \I__2029\ : Span12Mux_v
    port map (
            O => \N__9091\,
            I => \N__9088\
        );

    \I__2028\ : Odrv12
    port map (
            O => \N__9088\,
            I => \CLK40_PLL_i\
        );

    \I__2027\ : IoInMux
    port map (
            O => \N__9085\,
            I => \N__9082\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9082\,
            I => \N__9078\
        );

    \I__2025\ : IoInMux
    port map (
            O => \N__9081\,
            I => \N__9074\
        );

    \I__2024\ : Span4Mux_s2_v
    port map (
            O => \N__9078\,
            I => \N__9071\
        );

    \I__2023\ : IoInMux
    port map (
            O => \N__9077\,
            I => \N__9068\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__9074\,
            I => \N__9065\
        );

    \I__2021\ : Sp12to4
    port map (
            O => \N__9071\,
            I => \N__9062\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9068\,
            I => \N__9059\
        );

    \I__2019\ : Span4Mux_s3_h
    port map (
            O => \N__9065\,
            I => \N__9056\
        );

    \I__2018\ : Span12Mux_h
    port map (
            O => \N__9062\,
            I => \N__9053\
        );

    \I__2017\ : Span12Mux_s2_v
    port map (
            O => \N__9059\,
            I => \N__9050\
        );

    \I__2016\ : Span4Mux_h
    port map (
            O => \N__9056\,
            I => \N__9047\
        );

    \I__2015\ : Span12Mux_v
    port map (
            O => \N__9053\,
            I => \N__9042\
        );

    \I__2014\ : Span12Mux_v
    port map (
            O => \N__9050\,
            I => \N__9042\
        );

    \I__2013\ : Span4Mux_h
    port map (
            O => \N__9047\,
            I => \N__9039\
        );

    \I__2012\ : Span12Mux_h
    port map (
            O => \N__9042\,
            I => \N__9036\
        );

    \I__2011\ : Span4Mux_h
    port map (
            O => \N__9039\,
            I => \N__9033\
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9036\,
            I => \CLK40_PLL_i_i\
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__9033\,
            I => \CLK40_PLL_i_i\
        );

    \I__2008\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9024\
        );

    \I__2007\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9021\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9024\,
            I => \N__9018\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9021\,
            I => \N__9015\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__9018\,
            I => \N_334\
        );

    \I__2003\ : Odrv12
    port map (
            O => \N__9015\,
            I => \N_334\
        );

    \I__2002\ : InMux
    port map (
            O => \N__9010\,
            I => \N__9002\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__9009\,
            I => \N__8999\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__9008\,
            I => \N__8996\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9007\,
            I => \N__8991\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__9006\,
            I => \N__8988\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8985\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8982\
        );

    \I__1995\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8978\
        );

    \I__1994\ : InMux
    port map (
            O => \N__8996\,
            I => \N__8975\
        );

    \I__1993\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8972\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8965\
        );

    \I__1991\ : InMux
    port map (
            O => \N__8991\,
            I => \N__8965\
        );

    \I__1990\ : InMux
    port map (
            O => \N__8988\,
            I => \N__8960\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8985\,
            I => \N__8956\
        );

    \I__1988\ : Span4Mux_v
    port map (
            O => \N__8982\,
            I => \N__8953\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__8981\,
            I => \N__8950\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8945\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8975\,
            I => \N__8945\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8972\,
            I => \N__8942\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8939\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8936\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8965\,
            I => \N__8933\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8964\,
            I => \N__8928\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8963\,
            I => \N__8928\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__8960\,
            I => \N__8925\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8922\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__8956\,
            I => \N__8917\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__8953\,
            I => \N__8917\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8914\
        );

    \I__1973\ : Span4Mux_v
    port map (
            O => \N__8945\,
            I => \N__8901\
        );

    \I__1972\ : Span4Mux_v
    port map (
            O => \N__8942\,
            I => \N__8901\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N__8901\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N__8901\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__8933\,
            I => \N__8901\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8928\,
            I => \N__8901\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__8925\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8922\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1965\ : Odrv4
    port map (
            O => \N__8917\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8914\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1963\ : Odrv4
    port map (
            O => \N__8901\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1962\ : IoInMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__1960\ : Span4Mux_s1_v
    port map (
            O => \N__8884\,
            I => \N__8881\
        );

    \I__1959\ : Sp12to4
    port map (
            O => \N__8881\,
            I => \N__8878\
        );

    \I__1958\ : Span12Mux_h
    port map (
            O => \N__8878\,
            I => \N__8875\
        );

    \I__1957\ : Odrv12
    port map (
            O => \N__8875\,
            I => \ASn_c\
        );

    \I__1956\ : CEMux
    port map (
            O => \N__8872\,
            I => \N__8869\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8869\,
            I => \N__8866\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__8866\,
            I => \N__8863\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__8863\,
            I => \N__8860\
        );

    \I__1952\ : Odrv4
    port map (
            O => \N__8860\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__8857\,
            I => \N__8852\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8849\
        );

    \I__1949\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8846\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8841\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8827\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8827\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8824\
        );

    \I__1944\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8820\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8807\
        );

    \I__1942\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8800\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8800\
        );

    \I__1940\ : InMux
    port map (
            O => \N__8838\,
            I => \N__8800\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8797\
        );

    \I__1938\ : InMux
    port map (
            O => \N__8836\,
            I => \N__8790\
        );

    \I__1937\ : InMux
    port map (
            O => \N__8835\,
            I => \N__8790\
        );

    \I__1936\ : InMux
    port map (
            O => \N__8834\,
            I => \N__8790\
        );

    \I__1935\ : InMux
    port map (
            O => \N__8833\,
            I => \N__8787\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8832\,
            I => \N__8783\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__8827\,
            I => \N__8778\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__8824\,
            I => \N__8778\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8823\,
            I => \N__8775\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8820\,
            I => \N__8772\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8819\,
            I => \N__8765\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8818\,
            I => \N__8765\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8765\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8762\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8759\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8756\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8813\,
            I => \N__8753\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8812\,
            I => \N__8750\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8811\,
            I => \N__8747\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8810\,
            I => \N__8744\
        );

    \I__1919\ : Span4Mux_v
    port map (
            O => \N__8807\,
            I => \N__8738\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8800\,
            I => \N__8738\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8733\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8733\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8787\,
            I => \N__8730\
        );

    \I__1914\ : InMux
    port map (
            O => \N__8786\,
            I => \N__8727\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__8783\,
            I => \N__8720\
        );

    \I__1912\ : Span4Mux_v
    port map (
            O => \N__8778\,
            I => \N__8720\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__8775\,
            I => \N__8720\
        );

    \I__1910\ : Span4Mux_v
    port map (
            O => \N__8772\,
            I => \N__8709\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8709\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8709\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8759\,
            I => \N__8709\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8756\,
            I => \N__8709\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8753\,
            I => \N__8700\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8700\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8700\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8700\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__8743\,
            I => \N__8696\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__8738\,
            I => \N__8687\
        );

    \I__1899\ : Span4Mux_v
    port map (
            O => \N__8733\,
            I => \N__8687\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__8730\,
            I => \N__8687\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__8727\,
            I => \N__8682\
        );

    \I__1896\ : Sp12to4
    port map (
            O => \N__8720\,
            I => \N__8682\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__8709\,
            I => \N__8677\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__8700\,
            I => \N__8677\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8699\,
            I => \N__8668\
        );

    \I__1892\ : InMux
    port map (
            O => \N__8696\,
            I => \N__8668\
        );

    \I__1891\ : InMux
    port map (
            O => \N__8695\,
            I => \N__8668\
        );

    \I__1890\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8668\
        );

    \I__1889\ : Sp12to4
    port map (
            O => \N__8687\,
            I => \N__8663\
        );

    \I__1888\ : Span12Mux_v
    port map (
            O => \N__8682\,
            I => \N__8663\
        );

    \I__1887\ : Sp12to4
    port map (
            O => \N__8677\,
            I => \N__8658\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__8668\,
            I => \N__8658\
        );

    \I__1885\ : Span12Mux_h
    port map (
            O => \N__8663\,
            I => \N__8655\
        );

    \I__1884\ : Span12Mux_h
    port map (
            O => \N__8658\,
            I => \N__8652\
        );

    \I__1883\ : Odrv12
    port map (
            O => \N__8655\,
            I => \RESETn_c\
        );

    \I__1882\ : Odrv12
    port map (
            O => \N__8652\,
            I => \RESETn_c\
        );

    \I__1881\ : IoInMux
    port map (
            O => \N__8647\,
            I => \N__8644\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__8641\,
            I => \RESETn_c_i\
        );

    \I__1878\ : IoInMux
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8632\
        );

    \I__1876\ : Span4Mux_s3_v
    port map (
            O => \N__8632\,
            I => \N__8629\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__8629\,
            I => \N__8626\
        );

    \I__1874\ : Odrv4
    port map (
            O => \N__8626\,
            I => \N_353_i\
        );

    \I__1873\ : IoInMux
    port map (
            O => \N__8623\,
            I => \N__8620\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8620\,
            I => \N__8617\
        );

    \I__1871\ : Span4Mux_s2_v
    port map (
            O => \N__8617\,
            I => \N__8614\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__8614\,
            I => \N__8611\
        );

    \I__1869\ : Sp12to4
    port map (
            O => \N__8611\,
            I => \N__8608\
        );

    \I__1868\ : Odrv12
    port map (
            O => \N__8608\,
            I => \N_354_i\
        );

    \I__1867\ : IoInMux
    port map (
            O => \N__8605\,
            I => \N__8602\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__8602\,
            I => \N__8599\
        );

    \I__1865\ : IoSpan4Mux
    port map (
            O => \N__8599\,
            I => \N__8596\
        );

    \I__1864\ : Span4Mux_s3_v
    port map (
            O => \N__8596\,
            I => \N__8593\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8593\,
            I => \N_84_i\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8585\
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8589\,
            I => \N__8582\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__8588\,
            I => \N__8579\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8585\,
            I => \N__8576\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8573\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8570\
        );

    \I__1856\ : Span4Mux_v
    port map (
            O => \N__8576\,
            I => \N__8559\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__8573\,
            I => \N__8559\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8559\
        );

    \I__1853\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8556\
        );

    \I__1852\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8549\
        );

    \I__1851\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8549\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8549\
        );

    \I__1849\ : Span4Mux_h
    port map (
            O => \N__8559\,
            I => \N__8546\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8541\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__8549\,
            I => \N__8541\
        );

    \I__1846\ : Sp12to4
    port map (
            O => \N__8546\,
            I => \N__8538\
        );

    \I__1845\ : Span12Mux_v
    port map (
            O => \N__8541\,
            I => \N__8535\
        );

    \I__1844\ : Span12Mux_v
    port map (
            O => \N__8538\,
            I => \N__8532\
        );

    \I__1843\ : Span12Mux_h
    port map (
            O => \N__8535\,
            I => \N__8529\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8532\,
            I => \SIZ_c_0\
        );

    \I__1841\ : Odrv12
    port map (
            O => \N__8529\,
            I => \SIZ_c_0\
        );

    \I__1840\ : InMux
    port map (
            O => \N__8524\,
            I => \N__8521\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8521\,
            I => \N__8516\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8520\,
            I => \N__8513\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8506\
        );

    \I__1836\ : Span4Mux_h
    port map (
            O => \N__8516\,
            I => \N__8501\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8513\,
            I => \N__8501\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8512\,
            I => \N__8494\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8511\,
            I => \N__8494\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8510\,
            I => \N__8494\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8509\,
            I => \N__8491\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8506\,
            I => \N__8488\
        );

    \I__1829\ : Span4Mux_h
    port map (
            O => \N__8501\,
            I => \N__8485\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8478\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8491\,
            I => \N__8478\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__8488\,
            I => \N__8475\
        );

    \I__1825\ : Span4Mux_v
    port map (
            O => \N__8485\,
            I => \N__8472\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8484\,
            I => \N__8469\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8466\
        );

    \I__1822\ : Span12Mux_s10_v
    port map (
            O => \N__8478\,
            I => \N__8455\
        );

    \I__1821\ : Sp12to4
    port map (
            O => \N__8475\,
            I => \N__8455\
        );

    \I__1820\ : Sp12to4
    port map (
            O => \N__8472\,
            I => \N__8455\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8455\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8466\,
            I => \N__8455\
        );

    \I__1817\ : Span12Mux_h
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__8452\,
            I => \A_c_0\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8446\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__8446\,
            I => \N__8440\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8445\,
            I => \N__8437\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__8444\,
            I => \N__8434\
        );

    \I__1811\ : InMux
    port map (
            O => \N__8443\,
            I => \N__8430\
        );

    \I__1810\ : Span4Mux_v
    port map (
            O => \N__8440\,
            I => \N__8425\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8425\
        );

    \I__1808\ : InMux
    port map (
            O => \N__8434\,
            I => \N__8422\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8433\,
            I => \N__8418\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8430\,
            I => \N__8414\
        );

    \I__1805\ : Span4Mux_h
    port map (
            O => \N__8425\,
            I => \N__8409\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__8422\,
            I => \N__8409\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8402\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8402\
        );

    \I__1801\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8402\
        );

    \I__1800\ : Span4Mux_v
    port map (
            O => \N__8414\,
            I => \N__8399\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__8409\,
            I => \N__8393\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__8402\,
            I => \N__8393\
        );

    \I__1797\ : Span4Mux_v
    port map (
            O => \N__8399\,
            I => \N__8390\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8387\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__8393\,
            I => \N__8384\
        );

    \I__1794\ : Span4Mux_v
    port map (
            O => \N__8390\,
            I => \N__8381\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8387\,
            I => \N__8378\
        );

    \I__1792\ : Span4Mux_v
    port map (
            O => \N__8384\,
            I => \N__8375\
        );

    \I__1791\ : Sp12to4
    port map (
            O => \N__8381\,
            I => \N__8370\
        );

    \I__1790\ : Span12Mux_v
    port map (
            O => \N__8378\,
            I => \N__8370\
        );

    \I__1789\ : Span4Mux_h
    port map (
            O => \N__8375\,
            I => \N__8367\
        );

    \I__1788\ : Span12Mux_h
    port map (
            O => \N__8370\,
            I => \N__8364\
        );

    \I__1787\ : Sp12to4
    port map (
            O => \N__8367\,
            I => \N__8361\
        );

    \I__1786\ : Odrv12
    port map (
            O => \N__8364\,
            I => \SIZ_c_1\
        );

    \I__1785\ : Odrv12
    port map (
            O => \N__8361\,
            I => \SIZ_c_1\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__8356\,
            I => \N__8352\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8355\,
            I => \N__8349\
        );

    \I__1782\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8346\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__8349\,
            I => \N__8337\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__8346\,
            I => \N__8337\
        );

    \I__1779\ : CascadeMux
    port map (
            O => \N__8345\,
            I => \N__8334\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__8344\,
            I => \N__8330\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8325\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8325\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__8337\,
            I => \N__8322\
        );

    \I__1774\ : InMux
    port map (
            O => \N__8334\,
            I => \N__8315\
        );

    \I__1773\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8315\
        );

    \I__1772\ : InMux
    port map (
            O => \N__8330\,
            I => \N__8315\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__8325\,
            I => \N__8311\
        );

    \I__1770\ : Span4Mux_v
    port map (
            O => \N__8322\,
            I => \N__8308\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8315\,
            I => \N__8305\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8302\
        );

    \I__1767\ : Span12Mux_v
    port map (
            O => \N__8311\,
            I => \N__8295\
        );

    \I__1766\ : Sp12to4
    port map (
            O => \N__8308\,
            I => \N__8295\
        );

    \I__1765\ : Span12Mux_s7_v
    port map (
            O => \N__8305\,
            I => \N__8295\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8292\
        );

    \I__1763\ : Span12Mux_h
    port map (
            O => \N__8295\,
            I => \N__8289\
        );

    \I__1762\ : Span12Mux_h
    port map (
            O => \N__8292\,
            I => \N__8286\
        );

    \I__1761\ : Odrv12
    port map (
            O => \N__8289\,
            I => \A_c_1\
        );

    \I__1760\ : Odrv12
    port map (
            O => \N__8286\,
            I => \A_c_1\
        );

    \I__1759\ : IoInMux
    port map (
            O => \N__8281\,
            I => \N__8278\
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__8278\,
            I => \N__8275\
        );

    \I__1757\ : Span4Mux_s3_v
    port map (
            O => \N__8275\,
            I => \N__8272\
        );

    \I__1756\ : Span4Mux_h
    port map (
            O => \N__8272\,
            I => \N__8269\
        );

    \I__1755\ : Odrv4
    port map (
            O => \N__8269\,
            I => \N_355_i\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8263\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8263\,
            I => \N__8260\
        );

    \I__1752\ : Odrv4
    port map (
            O => \N__8260\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__8257\,
            I => \N__8249\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__8256\,
            I => \N__8246\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__8255\,
            I => \N__8242\
        );

    \I__1748\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8239\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__8253\,
            I => \N__8233\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__8252\,
            I => \N__8230\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8224\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8246\,
            I => \N__8219\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8219\
        );

    \I__1742\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8216\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8239\,
            I => \N__8213\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8238\,
            I => \N__8210\
        );

    \I__1739\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8207\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8202\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8233\,
            I => \N__8202\
        );

    \I__1736\ : InMux
    port map (
            O => \N__8230\,
            I => \N__8199\
        );

    \I__1735\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8194\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8194\
        );

    \I__1733\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8191\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__8224\,
            I => \N__8182\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8219\,
            I => \N__8175\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8216\,
            I => \N__8175\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__8213\,
            I => \N__8170\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8210\,
            I => \N__8170\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__8207\,
            I => \N__8165\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8165\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__8199\,
            I => \N__8158\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8194\,
            I => \N__8158\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8191\,
            I => \N__8158\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8150\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8150\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8141\
        );

    \I__1719\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8141\
        );

    \I__1718\ : InMux
    port map (
            O => \N__8186\,
            I => \N__8141\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8185\,
            I => \N__8141\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__8182\,
            I => \N__8138\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8181\,
            I => \N__8133\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8133\
        );

    \I__1713\ : Span4Mux_h
    port map (
            O => \N__8175\,
            I => \N__8124\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__8170\,
            I => \N__8124\
        );

    \I__1711\ : Span4Mux_v
    port map (
            O => \N__8165\,
            I => \N__8124\
        );

    \I__1710\ : Span4Mux_v
    port map (
            O => \N__8158\,
            I => \N__8124\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8121\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8156\,
            I => \N__8116\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8155\,
            I => \N__8116\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8150\,
            I => \N__8111\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__8141\,
            I => \N__8111\
        );

    \I__1704\ : Odrv4
    port map (
            O => \N__8138\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__8133\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1702\ : Odrv4
    port map (
            O => \N__8124\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8121\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8116\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__8111\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__8098\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\
        );

    \I__1697\ : IoInMux
    port map (
            O => \N__8095\,
            I => \N__8092\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__8092\,
            I => \N__8089\
        );

    \I__1695\ : IoSpan4Mux
    port map (
            O => \N__8089\,
            I => \N__8086\
        );

    \I__1694\ : Span4Mux_s3_v
    port map (
            O => \N__8086\,
            I => \N__8083\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__8083\,
            I => \N__8080\
        );

    \I__1692\ : Span4Mux_v
    port map (
            O => \N__8080\,
            I => \N__8077\
        );

    \I__1691\ : Span4Mux_v
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__8074\,
            I => \CMA_c_0\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8068\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8068\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1687\ : IoInMux
    port map (
            O => \N__8065\,
            I => \N__8062\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8062\,
            I => \N__8059\
        );

    \I__1685\ : IoSpan4Mux
    port map (
            O => \N__8059\,
            I => \N__8056\
        );

    \I__1684\ : Sp12to4
    port map (
            O => \N__8056\,
            I => \N__8053\
        );

    \I__1683\ : Span12Mux_s9_v
    port map (
            O => \N__8053\,
            I => \N__8050\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__8050\,
            I => \CMA_c_2\
        );

    \I__1681\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8037\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8037\
        );

    \I__1679\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8034\
        );

    \I__1678\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8029\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8029\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8026\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8037\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8034\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8029\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8026\,
            I => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__8017\,
            I => \N__8009\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8016\,
            I => \N__8005\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8015\,
            I => \N__7998\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8014\,
            I => \N__7998\
        );

    \I__1667\ : InMux
    port map (
            O => \N__8013\,
            I => \N__7998\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8012\,
            I => \N__7990\
        );

    \I__1665\ : InMux
    port map (
            O => \N__8009\,
            I => \N__7990\
        );

    \I__1664\ : InMux
    port map (
            O => \N__8008\,
            I => \N__7990\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__7985\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7998\,
            I => \N__7985\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__7997\,
            I => \N__7982\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7990\,
            I => \N__7977\
        );

    \I__1659\ : Span4Mux_h
    port map (
            O => \N__7985\,
            I => \N__7974\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7982\,
            I => \N__7967\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7981\,
            I => \N__7967\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7980\,
            I => \N__7967\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__7977\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__7974\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7967\,
            I => \U712_CHIP_RAM.N_337\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7957\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7957\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1650\ : IoInMux
    port map (
            O => \N__7954\,
            I => \N__7951\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7948\
        );

    \I__1648\ : IoSpan4Mux
    port map (
            O => \N__7948\,
            I => \N__7945\
        );

    \I__1647\ : Sp12to4
    port map (
            O => \N__7945\,
            I => \N__7942\
        );

    \I__1646\ : Span12Mux_s3_h
    port map (
            O => \N__7942\,
            I => \N__7939\
        );

    \I__1645\ : Span12Mux_h
    port map (
            O => \N__7939\,
            I => \N__7936\
        );

    \I__1644\ : Span12Mux_v
    port map (
            O => \N__7936\,
            I => \N__7933\
        );

    \I__1643\ : Odrv12
    port map (
            O => \N__7933\,
            I => \CMA_c_3\
        );

    \I__1642\ : CEMux
    port map (
            O => \N__7930\,
            I => \N__7927\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7927\,
            I => \N__7922\
        );

    \I__1640\ : CEMux
    port map (
            O => \N__7926\,
            I => \N__7919\
        );

    \I__1639\ : CEMux
    port map (
            O => \N__7925\,
            I => \N__7916\
        );

    \I__1638\ : Span4Mux_h
    port map (
            O => \N__7922\,
            I => \N__7908\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7919\,
            I => \N__7908\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7908\
        );

    \I__1635\ : CEMux
    port map (
            O => \N__7915\,
            I => \N__7905\
        );

    \I__1634\ : Span4Mux_v
    port map (
            O => \N__7908\,
            I => \N__7900\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7900\
        );

    \I__1632\ : Odrv4
    port map (
            O => \N__7900\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__7897\,
            I => \N__7894\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7891\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__7891\,
            I => \N__7888\
        );

    \I__1628\ : Span4Mux_h
    port map (
            O => \N__7888\,
            I => \N__7885\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__7885\,
            I => \U712_BYTE_ENABLE.N_441\
        );

    \I__1626\ : IoInMux
    port map (
            O => \N__7882\,
            I => \N__7879\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7879\,
            I => \N__7876\
        );

    \I__1624\ : IoSpan4Mux
    port map (
            O => \N__7876\,
            I => \N__7873\
        );

    \I__1623\ : Sp12to4
    port map (
            O => \N__7873\,
            I => \N__7870\
        );

    \I__1622\ : Span12Mux_s9_h
    port map (
            O => \N__7870\,
            I => \N__7867\
        );

    \I__1621\ : Span12Mux_v
    port map (
            O => \N__7867\,
            I => \N__7864\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__7864\,
            I => \N_34_i\
        );

    \I__1619\ : CascadeMux
    port map (
            O => \N__7861\,
            I => \U712_BYTE_ENABLE.N_451_cascade_\
        );

    \I__1618\ : IoInMux
    port map (
            O => \N__7858\,
            I => \N__7855\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7855\,
            I => \N__7852\
        );

    \I__1616\ : Span4Mux_s3_h
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__1615\ : Span4Mux_v
    port map (
            O => \N__7849\,
            I => \N__7846\
        );

    \I__1614\ : Sp12to4
    port map (
            O => \N__7846\,
            I => \N__7843\
        );

    \I__1613\ : Span12Mux_s11_h
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__1612\ : Span12Mux_v
    port map (
            O => \N__7840\,
            I => \N__7837\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__7837\,
            I => \N_200_i\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__7834\,
            I => \N__7828\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__7833\,
            I => \N__7825\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__7832\,
            I => \N__7822\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__7831\,
            I => \N__7813\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7828\,
            I => \N__7798\
        );

    \I__1605\ : InMux
    port map (
            O => \N__7825\,
            I => \N__7798\
        );

    \I__1604\ : InMux
    port map (
            O => \N__7822\,
            I => \N__7795\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7821\,
            I => \N__7792\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7820\,
            I => \N__7789\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7786\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7783\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7780\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7816\,
            I => \N__7777\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7773\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7812\,
            I => \N__7770\
        );

    \I__1595\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7767\
        );

    \I__1594\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7762\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7762\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__7808\,
            I => \N__7758\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7807\,
            I => \N__7749\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7806\,
            I => \N__7749\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7749\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7744\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7803\,
            I => \N__7744\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7798\,
            I => \N__7737\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7795\,
            I => \N__7737\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7792\,
            I => \N__7737\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7789\,
            I => \N__7734\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__7786\,
            I => \N__7731\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__7783\,
            I => \N__7728\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__7780\,
            I => \N__7725\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7777\,
            I => \N__7722\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7776\,
            I => \N__7719\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7773\,
            I => \N__7714\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7770\,
            I => \N__7714\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7767\,
            I => \N__7711\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7762\,
            I => \N__7708\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7705\
        );

    \I__1572\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7700\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7757\,
            I => \N__7700\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7756\,
            I => \N__7697\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7749\,
            I => \N__7694\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7744\,
            I => \N__7691\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__7737\,
            I => \N__7682\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__7734\,
            I => \N__7682\
        );

    \I__1565\ : Span4Mux_v
    port map (
            O => \N__7731\,
            I => \N__7682\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__7728\,
            I => \N__7682\
        );

    \I__1563\ : Odrv12
    port map (
            O => \N__7725\,
            I => \CPU_CYCLEm\
        );

    \I__1562\ : Odrv4
    port map (
            O => \N__7722\,
            I => \CPU_CYCLEm\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__7719\,
            I => \CPU_CYCLEm\
        );

    \I__1560\ : Odrv4
    port map (
            O => \N__7714\,
            I => \CPU_CYCLEm\
        );

    \I__1559\ : Odrv4
    port map (
            O => \N__7711\,
            I => \CPU_CYCLEm\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__7708\,
            I => \CPU_CYCLEm\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7705\,
            I => \CPU_CYCLEm\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__7700\,
            I => \CPU_CYCLEm\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__7697\,
            I => \CPU_CYCLEm\
        );

    \I__1554\ : Odrv4
    port map (
            O => \N__7694\,
            I => \CPU_CYCLEm\
        );

    \I__1553\ : Odrv12
    port map (
            O => \N__7691\,
            I => \CPU_CYCLEm\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__7682\,
            I => \CPU_CYCLEm\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7657\,
            I => \N__7651\
        );

    \I__1550\ : InMux
    port map (
            O => \N__7656\,
            I => \N__7646\
        );

    \I__1549\ : InMux
    port map (
            O => \N__7655\,
            I => \N__7646\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7643\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7651\,
            I => \N__7640\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__7646\,
            I => \N__7637\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7643\,
            I => \N__7634\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__7640\,
            I => \U712_BYTE_ENABLE.N_323_i\
        );

    \I__1543\ : Odrv4
    port map (
            O => \N__7637\,
            I => \U712_BYTE_ENABLE.N_323_i\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__7634\,
            I => \U712_BYTE_ENABLE.N_323_i\
        );

    \I__1541\ : CascadeMux
    port map (
            O => \N__7627\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\
        );

    \I__1540\ : IoInMux
    port map (
            O => \N__7624\,
            I => \N__7621\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7618\
        );

    \I__1538\ : IoSpan4Mux
    port map (
            O => \N__7618\,
            I => \N__7615\
        );

    \I__1537\ : Span4Mux_s3_h
    port map (
            O => \N__7615\,
            I => \N__7612\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__7612\,
            I => \N__7609\
        );

    \I__1535\ : Sp12to4
    port map (
            O => \N__7609\,
            I => \N__7606\
        );

    \I__1534\ : Span12Mux_h
    port map (
            O => \N__7606\,
            I => \N__7603\
        );

    \I__1533\ : Odrv12
    port map (
            O => \N__7603\,
            I => \CMA_c_4\
        );

    \I__1532\ : IoInMux
    port map (
            O => \N__7600\,
            I => \N__7597\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7597\,
            I => \N__7594\
        );

    \I__1530\ : Span12Mux_s5_v
    port map (
            O => \N__7594\,
            I => \N__7591\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7591\,
            I => \CMA_c_1\
        );

    \I__1528\ : IoInMux
    port map (
            O => \N__7588\,
            I => \N__7585\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7585\,
            I => \N__7582\
        );

    \I__1526\ : IoSpan4Mux
    port map (
            O => \N__7582\,
            I => \N__7579\
        );

    \I__1525\ : Sp12to4
    port map (
            O => \N__7579\,
            I => \N__7576\
        );

    \I__1524\ : Span12Mux_s7_v
    port map (
            O => \N__7576\,
            I => \N__7573\
        );

    \I__1523\ : Span12Mux_h
    port map (
            O => \N__7573\,
            I => \N__7570\
        );

    \I__1522\ : Odrv12
    port map (
            O => \N__7570\,
            I => \CMA_c_10\
        );

    \I__1521\ : IoInMux
    port map (
            O => \N__7567\,
            I => \N__7564\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__1519\ : IoSpan4Mux
    port map (
            O => \N__7561\,
            I => \N__7558\
        );

    \I__1518\ : Sp12to4
    port map (
            O => \N__7558\,
            I => \N__7555\
        );

    \I__1517\ : Span12Mux_s7_h
    port map (
            O => \N__7555\,
            I => \N__7552\
        );

    \I__1516\ : Span12Mux_v
    port map (
            O => \N__7552\,
            I => \N__7549\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__7549\,
            I => \CMA_c_6\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7543\
        );

    \I__1513\ : LocalMux
    port map (
            O => \N__7543\,
            I => \N__7540\
        );

    \I__1512\ : Odrv12
    port map (
            O => \N__7540\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1510\ : InMux
    port map (
            O => \N__7534\,
            I => \N__7531\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7531\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__7528\,
            I => \N__7525\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7525\,
            I => \N__7522\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__7522\,
            I => \N__7519\
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__7519\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1504\ : IoInMux
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7510\
        );

    \I__1502\ : IoSpan4Mux
    port map (
            O => \N__7510\,
            I => \N__7507\
        );

    \I__1501\ : Span4Mux_s2_v
    port map (
            O => \N__7507\,
            I => \N__7503\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7500\
        );

    \I__1499\ : Sp12to4
    port map (
            O => \N__7503\,
            I => \N__7497\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__7500\,
            I => \N__7494\
        );

    \I__1497\ : Span12Mux_s8_v
    port map (
            O => \N__7497\,
            I => \N__7491\
        );

    \I__1496\ : Span4Mux_v
    port map (
            O => \N__7494\,
            I => \N__7488\
        );

    \I__1495\ : Span12Mux_v
    port map (
            O => \N__7491\,
            I => \N__7483\
        );

    \I__1494\ : Sp12to4
    port map (
            O => \N__7488\,
            I => \N__7483\
        );

    \I__1493\ : Span12Mux_h
    port map (
            O => \N__7483\,
            I => \N__7480\
        );

    \I__1492\ : Odrv12
    port map (
            O => \N__7480\,
            I => \A_c_10\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7474\,
            I => \U712_CHIP_RAM.N_382\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7468\,
            I => \N__7465\
        );

    \I__1487\ : Span4Mux_h
    port map (
            O => \N__7465\,
            I => \N__7462\
        );

    \I__1486\ : Sp12to4
    port map (
            O => \N__7462\,
            I => \N__7459\
        );

    \I__1485\ : Span12Mux_v
    port map (
            O => \N__7459\,
            I => \N__7456\
        );

    \I__1484\ : Span12Mux_h
    port map (
            O => \N__7456\,
            I => \N__7453\
        );

    \I__1483\ : Odrv12
    port map (
            O => \N__7453\,
            I => \A_c_3\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7450\,
            I => \N__7447\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7447\,
            I => \U712_CHIP_RAM.N_374\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__7444\,
            I => \N__7441\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7438\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7438\,
            I => \N__7435\
        );

    \I__1477\ : Span4Mux_h
    port map (
            O => \N__7435\,
            I => \N__7432\
        );

    \I__1476\ : Odrv4
    port map (
            O => \N__7432\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7429\,
            I => \N__7424\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7421\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7418\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__7424\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7421\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7418\,
            I => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\
        );

    \I__1469\ : IoInMux
    port map (
            O => \N__7411\,
            I => \N__7408\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7405\
        );

    \I__1467\ : IoSpan4Mux
    port map (
            O => \N__7405\,
            I => \N__7402\
        );

    \I__1466\ : Span4Mux_s2_v
    port map (
            O => \N__7402\,
            I => \N__7399\
        );

    \I__1465\ : Sp12to4
    port map (
            O => \N__7399\,
            I => \N__7396\
        );

    \I__1464\ : Span12Mux_h
    port map (
            O => \N__7396\,
            I => \N__7392\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7395\,
            I => \N__7389\
        );

    \I__1462\ : Odrv12
    port map (
            O => \N__7392\,
            I => \LDSn_c\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7389\,
            I => \LDSn_c\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7384\,
            I => \N__7381\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7381\,
            I => \U712_REG_SM.N_446\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__7378\,
            I => \N__7375\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7372\
        );

    \I__1456\ : IoSpan4Mux
    port map (
            O => \N__7372\,
            I => \N__7369\
        );

    \I__1455\ : Span4Mux_s3_v
    port map (
            O => \N__7369\,
            I => \N__7366\
        );

    \I__1454\ : Span4Mux_v
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7363\,
            I => \N_435\
        );

    \I__1452\ : IoInMux
    port map (
            O => \N__7360\,
            I => \N__7357\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7354\
        );

    \I__1450\ : Span4Mux_s2_v
    port map (
            O => \N__7354\,
            I => \N__7351\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__7351\,
            I => \N__7348\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__7348\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1447\ : IoInMux
    port map (
            O => \N__7345\,
            I => \N__7342\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7342\,
            I => \N__7339\
        );

    \I__1445\ : Span12Mux_s2_v
    port map (
            O => \N__7339\,
            I => \N__7336\
        );

    \I__1444\ : Span12Mux_h
    port map (
            O => \N__7336\,
            I => \N__7333\
        );

    \I__1443\ : Odrv12
    port map (
            O => \N__7333\,
            I => \CASn_c\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \N__7325\
        );

    \I__1441\ : InMux
    port map (
            O => \N__7329\,
            I => \N__7320\
        );

    \I__1440\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7320\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7325\,
            I => \N__7317\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__7320\,
            I => \N__7312\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7317\,
            I => \N__7312\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__7312\,
            I => \N__7308\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7305\
        );

    \I__1434\ : Span4Mux_h
    port map (
            O => \N__7308\,
            I => \N__7298\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__7305\,
            I => \N__7298\
        );

    \I__1432\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7295\
        );

    \I__1431\ : InMux
    port map (
            O => \N__7303\,
            I => \N__7292\
        );

    \I__1430\ : Odrv4
    port map (
            O => \N__7298\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__7295\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7292\,
            I => \U712_CHIP_RAM.N_340\
        );

    \I__1427\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7281\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__7284\,
            I => \N__7273\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7281\,
            I => \N__7267\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7280\,
            I => \N__7262\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7279\,
            I => \N__7262\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__7278\,
            I => \N__7259\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7277\,
            I => \N__7255\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7276\,
            I => \N__7249\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7244\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7244\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7271\,
            I => \N__7239\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7270\,
            I => \N__7239\
        );

    \I__1415\ : Span4Mux_h
    port map (
            O => \N__7267\,
            I => \N__7234\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__7262\,
            I => \N__7234\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7231\
        );

    \I__1412\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7228\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7255\,
            I => \N__7225\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7220\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7253\,
            I => \N__7220\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7217\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__7249\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__7244\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1405\ : LocalMux
    port map (
            O => \N__7239\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1404\ : Odrv4
    port map (
            O => \N__7234\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7231\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7228\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1401\ : Odrv12
    port map (
            O => \N__7225\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__7220\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7217\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7194\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7197\,
            I => \N__7187\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7194\,
            I => \N__7182\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7179\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__7192\,
            I => \N__7173\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__7191\,
            I => \N__7170\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7190\,
            I => \N__7166\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7187\,
            I => \N__7163\
        );

    \I__1390\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7158\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7158\
        );

    \I__1388\ : Span4Mux_h
    port map (
            O => \N__7182\,
            I => \N__7149\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__7179\,
            I => \N__7146\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7143\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7140\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7137\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7130\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7170\,
            I => \N__7130\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7169\,
            I => \N__7130\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7166\,
            I => \N__7123\
        );

    \I__1379\ : Span4Mux_h
    port map (
            O => \N__7163\,
            I => \N__7123\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__7158\,
            I => \N__7123\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7157\,
            I => \N__7118\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7156\,
            I => \N__7118\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7155\,
            I => \N__7111\
        );

    \I__1374\ : InMux
    port map (
            O => \N__7154\,
            I => \N__7111\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7111\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7108\
        );

    \I__1371\ : Odrv4
    port map (
            O => \N__7149\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__7146\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7143\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7140\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__7137\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7130\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1365\ : Odrv4
    port map (
            O => \N__7123\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7118\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7111\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7108\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7084\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7084\,
            I => \N__7081\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__7081\,
            I => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7075\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__7066\,
            I => \U712_CHIP_RAM.DBENn_8_0\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1351\ : Odrv12
    port map (
            O => \N__7057\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1350\ : IoInMux
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1348\ : Span12Mux_s5_h
    port map (
            O => \N__7048\,
            I => \N__7045\
        );

    \I__1347\ : Span12Mux_v
    port map (
            O => \N__7045\,
            I => \N__7042\
        );

    \I__1346\ : Odrv12
    port map (
            O => \N__7042\,
            I => \CMA_c_5\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7036\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__7036\,
            I => \N__7033\
        );

    \I__1343\ : Odrv12
    port map (
            O => \N__7033\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1342\ : IoInMux
    port map (
            O => \N__7030\,
            I => \N__7027\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7027\,
            I => \N__7024\
        );

    \I__1340\ : IoSpan4Mux
    port map (
            O => \N__7024\,
            I => \N__7021\
        );

    \I__1339\ : Sp12to4
    port map (
            O => \N__7021\,
            I => \N__7018\
        );

    \I__1338\ : Span12Mux_s7_h
    port map (
            O => \N__7018\,
            I => \N__7015\
        );

    \I__1337\ : Span12Mux_v
    port map (
            O => \N__7015\,
            I => \N__7012\
        );

    \I__1336\ : Odrv12
    port map (
            O => \N__7012\,
            I => \CMA_c_7\
        );

    \I__1335\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \U712_BYTE_ENABLE.N_443_cascade_\
        );

    \I__1334\ : IoInMux
    port map (
            O => \N__7006\,
            I => \N__7003\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7003\,
            I => \N__7000\
        );

    \I__1332\ : IoSpan4Mux
    port map (
            O => \N__7000\,
            I => \N__6997\
        );

    \I__1331\ : IoSpan4Mux
    port map (
            O => \N__6997\,
            I => \N__6994\
        );

    \I__1330\ : Sp12to4
    port map (
            O => \N__6994\,
            I => \N__6991\
        );

    \I__1329\ : Span12Mux_s7_v
    port map (
            O => \N__6991\,
            I => \N__6988\
        );

    \I__1328\ : Span12Mux_h
    port map (
            O => \N__6988\,
            I => \N__6985\
        );

    \I__1327\ : Odrv12
    port map (
            O => \N__6985\,
            I => \N_32_i\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6979\,
            I => \N__6976\
        );

    \I__1324\ : Span4Mux_h
    port map (
            O => \N__6976\,
            I => \N__6973\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__6973\,
            I => \N__6970\
        );

    \I__1322\ : Sp12to4
    port map (
            O => \N__6970\,
            I => \N__6967\
        );

    \I__1321\ : Span12Mux_h
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__1320\ : Odrv12
    port map (
            O => \N__6964\,
            I => \A_c_20\
        );

    \I__1319\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6958\,
            I => \N__6955\
        );

    \I__1317\ : Odrv12
    port map (
            O => \N__6955\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6946\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6943\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6940\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6949\,
            I => \N__6937\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__6946\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6943\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6940\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6937\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_2\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6924\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6921\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6924\,
            I => \U712_REG_SM.N_348\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6921\,
            I => \U712_REG_SM.N_348\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__6916\,
            I => \U712_REG_SM.N_462_cascade_\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6910\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6910\,
            I => \U712_REG_SM.N_399\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6907\,
            I => \N__6901\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6901\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__6901\,
            I => \N__6898\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__6898\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__6895\,
            I => \U712_CHIP_RAM.N_440_cascade_\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6892\,
            I => \N__6889\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6889\,
            I => \U712_CHIP_RAM.N_439\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\
        );

    \I__1293\ : CEMux
    port map (
            O => \N__6883\,
            I => \N__6880\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6880\,
            I => \N__6877\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__6877\,
            I => \N__6874\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__6874\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__6871\,
            I => \N__6866\
        );

    \I__1288\ : InMux
    port map (
            O => \N__6870\,
            I => \N__6862\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6869\,
            I => \N__6856\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6866\,
            I => \N__6856\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__6865\,
            I => \N__6845\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__6862\,
            I => \N__6842\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6861\,
            I => \N__6839\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6856\,
            I => \N__6836\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__6855\,
            I => \N__6833\
        );

    \I__1280\ : CascadeMux
    port map (
            O => \N__6854\,
            I => \N__6828\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6853\,
            I => \N__6825\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6852\,
            I => \N__6818\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6818\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6818\
        );

    \I__1275\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6815\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6848\,
            I => \N__6812\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6845\,
            I => \N__6809\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__6842\,
            I => \N__6804\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6839\,
            I => \N__6804\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__6836\,
            I => \N__6801\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6798\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6832\,
            I => \N__6791\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6831\,
            I => \N__6791\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6791\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6825\,
            I => \N__6786\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6818\,
            I => \N__6786\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6815\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6812\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6809\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__6804\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__6801\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6798\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6791\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__6786\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1255\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6766\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6766\,
            I => \N__6763\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__6763\,
            I => \N__6758\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6755\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6752\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__6758\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6755\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6752\,
            I => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6742\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6742\,
            I => \U712_CHIP_RAM.N_507\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__6739\,
            I => \N__6732\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__6738\,
            I => \N__6728\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6721\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6721\
        );

    \I__1241\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6718\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6732\,
            I => \N__6715\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6710\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6710\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6727\,
            I => \N__6707\
        );

    \I__1236\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6704\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6701\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__6718\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6715\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__6710\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__6707\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__6704\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__6701\,
            I => \U712_CHIP_RAM.N_504\
        );

    \I__1228\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6684\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6681\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6684\,
            I => \N__6678\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6681\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__6678\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\
        );

    \I__1223\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6667\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__6667\,
            I => \U712_CHIP_RAM.N_48\
        );

    \I__1220\ : IoInMux
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1218\ : IoSpan4Mux
    port map (
            O => \N__6658\,
            I => \N__6655\
        );

    \I__1217\ : IoSpan4Mux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1216\ : Span4Mux_s3_v
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1215\ : Sp12to4
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1214\ : Span12Mux_s11_v
    port map (
            O => \N__6646\,
            I => \N__6642\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6645\,
            I => \N__6639\
        );

    \I__1212\ : Odrv12
    port map (
            O => \N__6642\,
            I => \LATCH_CLK_c\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__6639\,
            I => \LATCH_CLK_c\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6631\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__6628\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6625\,
            I => \N__6622\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6622\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6615\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6612\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6615\,
            I => \N__6608\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__6612\,
            I => \N__6605\
        );

    \I__1201\ : InMux
    port map (
            O => \N__6611\,
            I => \N__6602\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__6608\,
            I => \N__6597\
        );

    \I__1199\ : Span4Mux_h
    port map (
            O => \N__6605\,
            I => \N__6594\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6591\
        );

    \I__1197\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6588\
        );

    \I__1196\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6585\
        );

    \I__1195\ : Odrv4
    port map (
            O => \N__6597\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__6594\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1193\ : Odrv4
    port map (
            O => \N__6591\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6588\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6585\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6574\,
            I => \N__6571\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6566\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6570\,
            I => \N__6563\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6560\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__6566\,
            I => \N__6557\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6563\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__6560\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1183\ : Odrv4
    port map (
            O => \N__6557\,
            I => \U712_CHIP_RAM.N_327\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__6550\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\
        );

    \I__1181\ : InMux
    port map (
            O => \N__6547\,
            I => \N__6544\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6544\,
            I => \U712_CHIP_RAM.N_433\
        );

    \I__1179\ : InMux
    port map (
            O => \N__6541\,
            I => \N__6532\
        );

    \I__1178\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6529\
        );

    \I__1177\ : CascadeMux
    port map (
            O => \N__6539\,
            I => \N__6526\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__6538\,
            I => \N__6523\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6519\
        );

    \I__1174\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6516\
        );

    \I__1173\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6513\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6532\,
            I => \N__6508\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6529\,
            I => \N__6508\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6503\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6503\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6500\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__6519\,
            I => \N__6497\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6516\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1164\ : Odrv4
    port map (
            O => \N__6508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6503\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__6497\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6481\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__6481\,
            I => \N__6476\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6480\,
            I => \N__6473\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6479\,
            I => \N__6470\
        );

    \I__1156\ : Span4Mux_h
    port map (
            O => \N__6476\,
            I => \N__6467\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6473\,
            I => \N__6464\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6470\,
            I => \U712_CHIP_RAM.N_499\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__6467\,
            I => \U712_CHIP_RAM.N_499\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__6464\,
            I => \U712_CHIP_RAM.N_499\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6457\,
            I => \U712_CHIP_RAM.N_499_cascade_\
        );

    \I__1150\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6447\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6453\,
            I => \N__6447\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6444\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6441\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6444\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__1145\ : Odrv4
    port map (
            O => \N__6441\,
            I => \U712_CHIP_RAM.N_341\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__6436\,
            I => \U712_CHIP_RAM.N_507_cascade_\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__6430\,
            I => \U712_CHIP_RAM.N_438\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__6427\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6418\
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__6418\,
            I => \N__6413\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6417\,
            I => \N__6408\
        );

    \I__1136\ : InMux
    port map (
            O => \N__6416\,
            I => \N__6408\
        );

    \I__1135\ : Span4Mux_h
    port map (
            O => \N__6413\,
            I => \N__6399\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6408\,
            I => \N__6399\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__6407\,
            I => \N__6394\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__6406\,
            I => \N__6388\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6405\,
            I => \N__6385\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6382\
        );

    \I__1129\ : Sp12to4
    port map (
            O => \N__6399\,
            I => \N__6379\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6398\,
            I => \N__6376\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6367\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6394\,
            I => \N__6367\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6393\,
            I => \N__6367\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6367\
        );

    \I__1123\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6362\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6362\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6385\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__6382\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1119\ : Odrv12
    port map (
            O => \N__6379\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__6376\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6367\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6362\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1115\ : IoInMux
    port map (
            O => \N__6349\,
            I => \N__6346\
        );

    \I__1114\ : LocalMux
    port map (
            O => \N__6346\,
            I => \N__6343\
        );

    \I__1113\ : Span4Mux_s3_v
    port map (
            O => \N__6343\,
            I => \N__6340\
        );

    \I__1112\ : Sp12to4
    port map (
            O => \N__6340\,
            I => \N__6337\
        );

    \I__1111\ : Span12Mux_h
    port map (
            O => \N__6337\,
            I => \N__6333\
        );

    \I__1110\ : InMux
    port map (
            O => \N__6336\,
            I => \N__6330\
        );

    \I__1109\ : Odrv12
    port map (
            O => \N__6333\,
            I => \UDSn_c\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6330\,
            I => \UDSn_c\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6322\,
            I => \U712_REG_SM.N_447\
        );

    \I__1105\ : IoInMux
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1103\ : Span12Mux_s10_v
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1102\ : Odrv12
    port map (
            O => \N__6310\,
            I => \RASn_c\
        );

    \I__1101\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6304\,
            I => \N__6301\
        );

    \I__1099\ : Span4Mux_h
    port map (
            O => \N__6301\,
            I => \N__6298\
        );

    \I__1098\ : Sp12to4
    port map (
            O => \N__6298\,
            I => \N__6295\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6292\,
            I => \A_c_19\
        );

    \I__1095\ : IoInMux
    port map (
            O => \N__6289\,
            I => \N__6286\
        );

    \I__1094\ : LocalMux
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__1093\ : IoSpan4Mux
    port map (
            O => \N__6283\,
            I => \N__6280\
        );

    \I__1092\ : IoSpan4Mux
    port map (
            O => \N__6280\,
            I => \N__6277\
        );

    \I__1091\ : Span4Mux_s2_h
    port map (
            O => \N__6277\,
            I => \N__6274\
        );

    \I__1090\ : Sp12to4
    port map (
            O => \N__6274\,
            I => \N__6271\
        );

    \I__1089\ : Span12Mux_s9_h
    port map (
            O => \N__6271\,
            I => \N__6268\
        );

    \I__1088\ : Odrv12
    port map (
            O => \N__6268\,
            I => \CMA_c_9\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6262\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6257\
        );

    \I__1085\ : InMux
    port map (
            O => \N__6261\,
            I => \N__6254\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6251\
        );

    \I__1083\ : Span4Mux_v
    port map (
            O => \N__6257\,
            I => \N__6243\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6243\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__6251\,
            I => \N__6240\
        );

    \I__1080\ : InMux
    port map (
            O => \N__6250\,
            I => \N__6235\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6235\
        );

    \I__1078\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6232\
        );

    \I__1077\ : Span4Mux_h
    port map (
            O => \N__6243\,
            I => \N__6227\
        );

    \I__1076\ : Span4Mux_h
    port map (
            O => \N__6240\,
            I => \N__6227\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6224\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__6232\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1073\ : Odrv4
    port map (
            O => \N__6227\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1072\ : Odrv4
    port map (
            O => \N__6224\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6214\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6214\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6208\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6208\,
            I => \N__6205\
        );

    \I__1067\ : Span4Mux_v
    port map (
            O => \N__6205\,
            I => \N__6202\
        );

    \I__1066\ : Span4Mux_v
    port map (
            O => \N__6202\,
            I => \N__6199\
        );

    \I__1065\ : Sp12to4
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1064\ : Span12Mux_h
    port map (
            O => \N__6196\,
            I => \N__6193\
        );

    \I__1063\ : Odrv12
    port map (
            O => \N__6193\,
            I => \A_c_17\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6190\,
            I => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\
        );

    \I__1061\ : IoInMux
    port map (
            O => \N__6187\,
            I => \N__6184\
        );

    \I__1060\ : LocalMux
    port map (
            O => \N__6184\,
            I => \N__6181\
        );

    \I__1059\ : IoSpan4Mux
    port map (
            O => \N__6181\,
            I => \N__6178\
        );

    \I__1058\ : Span4Mux_s2_h
    port map (
            O => \N__6178\,
            I => \N__6175\
        );

    \I__1057\ : Span4Mux_h
    port map (
            O => \N__6175\,
            I => \N__6172\
        );

    \I__1056\ : Sp12to4
    port map (
            O => \N__6172\,
            I => \N__6169\
        );

    \I__1055\ : Span12Mux_h
    port map (
            O => \N__6169\,
            I => \N__6166\
        );

    \I__1054\ : Odrv12
    port map (
            O => \N__6166\,
            I => \CMA_c_8\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__6163\,
            I => \N__6160\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6157\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6157\,
            I => \N__6154\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__6154\,
            I => \N__6151\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6151\,
            I => \U712_CHIP_RAM.N_432\
        );

    \I__1048\ : IoInMux
    port map (
            O => \N__6148\,
            I => \N__6145\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1046\ : IoSpan4Mux
    port map (
            O => \N__6142\,
            I => \N__6139\
        );

    \I__1045\ : Span4Mux_s1_v
    port map (
            O => \N__6139\,
            I => \N__6136\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__6136\,
            I => \N__6133\
        );

    \I__1043\ : Span4Mux_v
    port map (
            O => \N__6133\,
            I => \N__6129\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6132\,
            I => \N__6126\
        );

    \I__1041\ : Odrv4
    port map (
            O => \N__6129\,
            I => \BANK0_c\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6126\,
            I => \BANK0_c\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6121\,
            I => \N__6118\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6118\,
            I => \N__6114\
        );

    \I__1037\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6111\
        );

    \I__1036\ : Odrv12
    port map (
            O => \N__6114\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6111\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__1034\ : CascadeMux
    port map (
            O => \N__6106\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_4_cascade_\
        );

    \I__1033\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6100\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6100\,
            I => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6093\
        );

    \I__1030\ : CascadeMux
    port map (
            O => \N__6096\,
            I => \N__6090\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6093\,
            I => \N__6087\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6090\,
            I => \N__6084\
        );

    \I__1027\ : Span4Mux_h
    port map (
            O => \N__6087\,
            I => \N__6080\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6077\
        );

    \I__1025\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6074\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6080\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1023\ : Odrv4
    port map (
            O => \N__6077\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6074\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6064\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6064\,
            I => \U712_REG_SM.STATE_COUNTc_0_0\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__6061\,
            I => \U712_REG_SM.N_348_cascade_\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6054\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6057\,
            I => \N__6051\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__6054\,
            I => \U712_REG_SM.N_347\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6051\,
            I => \U712_REG_SM.N_347\
        );

    \I__1014\ : CascadeMux
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6035\
        );

    \I__1012\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6035\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6043\,
            I => \N__6032\
        );

    \I__1010\ : InMux
    port map (
            O => \N__6040\,
            I => \N__6029\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__6035\,
            I => \N__6024\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6024\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__6029\,
            I => \REG_TACK\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__6024\,
            I => \REG_TACK\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6019\,
            I => \N__6014\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__6018\,
            I => \N__6011\
        );

    \I__1003\ : InMux
    port map (
            O => \N__6017\,
            I => \N__6005\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__6014\,
            I => \N__6002\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6011\,
            I => \N__5999\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6010\,
            I => \N__5996\
        );

    \I__999\ : InMux
    port map (
            O => \N__6009\,
            I => \N__5993\
        );

    \I__998\ : InMux
    port map (
            O => \N__6008\,
            I => \N__5990\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__6005\,
            I => \N__5987\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__6002\,
            I => \N__5982\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5999\,
            I => \N__5982\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5996\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5993\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5990\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__991\ : Odrv4
    port map (
            O => \N__5987\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__990\ : Odrv4
    port map (
            O => \N__5982\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_1\
        );

    \I__989\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5962\
        );

    \I__988\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5962\
        );

    \I__987\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5959\
        );

    \I__986\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5954\
        );

    \I__985\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5954\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5962\,
            I => \N__5951\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5959\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5954\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__981\ : Odrv4
    port map (
            O => \N__5951\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_4\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__5944\,
            I => \U712_REG_SM.N_399_cascade_\
        );

    \I__979\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5937\
        );

    \I__978\ : InMux
    port map (
            O => \N__5940\,
            I => \N__5934\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5937\,
            I => \N__5931\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__5934\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__975\ : Odrv12
    port map (
            O => \N__5931\,
            I => \U712_REG_SM.WRITE_CYCLEZ0\
        );

    \I__974\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5923\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__5923\,
            I => \U712_REG_SM.N_212\
        );

    \I__972\ : InMux
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__5919\,
            I => \N__5911\
        );

    \I__970\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5903\
        );

    \I__969\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5903\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5898\
        );

    \I__967\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5894\
        );

    \I__966\ : InMux
    port map (
            O => \N__5910\,
            I => \N__5891\
        );

    \I__965\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5886\
        );

    \I__964\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5886\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5903\,
            I => \N__5883\
        );

    \I__962\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5880\
        );

    \I__961\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5877\
        );

    \I__960\ : Span4Mux_h
    port map (
            O => \N__5898\,
            I => \N__5874\
        );

    \I__959\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5871\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5894\,
            I => \N__5868\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5859\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5886\,
            I => \N__5859\
        );

    \I__955\ : Span4Mux_v
    port map (
            O => \N__5883\,
            I => \N__5859\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5880\,
            I => \N__5859\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__5877\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__5874\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5871\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__950\ : Odrv4
    port map (
            O => \N__5868\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__949\ : Odrv4
    port map (
            O => \N__5859\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__5848\,
            I => \N__5842\
        );

    \I__947\ : InMux
    port map (
            O => \N__5847\,
            I => \N__5837\
        );

    \I__946\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5832\
        );

    \I__945\ : InMux
    port map (
            O => \N__5845\,
            I => \N__5832\
        );

    \I__944\ : InMux
    port map (
            O => \N__5842\,
            I => \N__5829\
        );

    \I__943\ : InMux
    port map (
            O => \N__5841\,
            I => \N__5826\
        );

    \I__942\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5823\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__5837\,
            I => \N__5818\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5832\,
            I => \N__5818\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5829\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5826\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5823\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__936\ : Odrv4
    port map (
            O => \N__5818\,
            I => \U712_REG_SM.STATE_COUNTZ0Z_3\
        );

    \I__935\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__5806\,
            I => \U712_REG_SM.N_458\
        );

    \I__933\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5797\
        );

    \I__932\ : InMux
    port map (
            O => \N__5802\,
            I => \N__5792\
        );

    \I__931\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5792\
        );

    \I__930\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5789\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5797\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5792\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5789\,
            I => \U712_CHIP_RAM.N_508\
        );

    \I__926\ : InMux
    port map (
            O => \N__5782\,
            I => \N__5778\
        );

    \I__925\ : InMux
    port map (
            O => \N__5781\,
            I => \N__5775\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5772\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U712_CHIP_RAM.N_610\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__5772\,
            I => \U712_CHIP_RAM.N_610\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__920\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5760\
        );

    \I__919\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5757\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5751\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5751\
        );

    \I__916\ : InMux
    port map (
            O => \N__5756\,
            I => \N__5748\
        );

    \I__915\ : Odrv4
    port map (
            O => \N__5751\,
            I => \U712_CHIP_RAM.N_608\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5748\,
            I => \U712_CHIP_RAM.N_608\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__5743\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\
        );

    \I__912\ : InMux
    port map (
            O => \N__5740\,
            I => \N__5737\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__5737\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_2\
        );

    \I__910\ : InMux
    port map (
            O => \N__5734\,
            I => \N__5731\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5731\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\
        );

    \I__908\ : InMux
    port map (
            O => \N__5728\,
            I => \N__5725\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5725\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\
        );

    \I__906\ : InMux
    port map (
            O => \N__5722\,
            I => \N__5718\
        );

    \I__905\ : InMux
    port map (
            O => \N__5721\,
            I => \N__5715\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5718\,
            I => \N__5712\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5709\
        );

    \I__902\ : Span4Mux_v
    port map (
            O => \N__5712\,
            I => \N__5706\
        );

    \I__901\ : Span4Mux_v
    port map (
            O => \N__5709\,
            I => \N__5703\
        );

    \I__900\ : Span4Mux_h
    port map (
            O => \N__5706\,
            I => \N__5700\
        );

    \I__899\ : Sp12to4
    port map (
            O => \N__5703\,
            I => \N__5697\
        );

    \I__898\ : Sp12to4
    port map (
            O => \N__5700\,
            I => \N__5692\
        );

    \I__897\ : Span12Mux_h
    port map (
            O => \N__5697\,
            I => \N__5692\
        );

    \I__896\ : Span12Mux_v
    port map (
            O => \N__5692\,
            I => \N__5689\
        );

    \I__895\ : Odrv12
    port map (
            O => \N__5689\,
            I => \AWEn_c\
        );

    \I__894\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5683\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5683\,
            I => \U712_CHIP_RAM.N_361\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__891\ : InMux
    port map (
            O => \N__5677\,
            I => \N__5670\
        );

    \I__890\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5670\
        );

    \I__889\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5667\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5670\,
            I => \N__5664\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5667\,
            I => \N__5661\
        );

    \I__886\ : Span4Mux_v
    port map (
            O => \N__5664\,
            I => \N__5658\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__5661\,
            I => \N__5655\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__5658\,
            I => \CPU_TACKm\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__5655\,
            I => \CPU_TACKm\
        );

    \I__882\ : InMux
    port map (
            O => \N__5650\,
            I => \N__5643\
        );

    \I__881\ : InMux
    port map (
            O => \N__5649\,
            I => \N__5643\
        );

    \I__880\ : InMux
    port map (
            O => \N__5648\,
            I => \N__5640\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__5643\,
            I => \N__5635\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__5640\,
            I => \N__5635\
        );

    \I__877\ : Odrv4
    port map (
            O => \N__5635\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__876\ : InMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5626\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__5626\,
            I => \U712_CYCLE_TERM.N_350\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__5623\,
            I => \N__5620\
        );

    \I__872\ : InMux
    port map (
            O => \N__5620\,
            I => \N__5617\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5614\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\
        );

    \I__869\ : CascadeMux
    port map (
            O => \N__5611\,
            I => \N__5608\
        );

    \I__868\ : InMux
    port map (
            O => \N__5608\,
            I => \N__5605\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5605\,
            I => \N__5600\
        );

    \I__866\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5597\
        );

    \I__865\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5593\
        );

    \I__864\ : Span4Mux_h
    port map (
            O => \N__5600\,
            I => \N__5590\
        );

    \I__863\ : LocalMux
    port map (
            O => \N__5597\,
            I => \N__5587\
        );

    \I__862\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5584\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__5593\,
            I => \U712_CHIP_RAM.N_515\
        );

    \I__860\ : Odrv4
    port map (
            O => \N__5590\,
            I => \U712_CHIP_RAM.N_515\
        );

    \I__859\ : Odrv4
    port map (
            O => \N__5587\,
            I => \U712_CHIP_RAM.N_515\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5584\,
            I => \U712_CHIP_RAM.N_515\
        );

    \I__857\ : InMux
    port map (
            O => \N__5575\,
            I => \N__5571\
        );

    \I__856\ : InMux
    port map (
            O => \N__5574\,
            I => \N__5568\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5571\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5568\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__853\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5559\
        );

    \I__852\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5556\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5559\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5556\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__849\ : InMux
    port map (
            O => \N__5551\,
            I => \N__5547\
        );

    \I__848\ : InMux
    port map (
            O => \N__5550\,
            I => \N__5544\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5547\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5544\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__845\ : CascadeMux
    port map (
            O => \N__5539\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7_cascade_\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__5536\,
            I => \U712_CHIP_RAM.N_504_cascade_\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__5533\,
            I => \U712_CHIP_RAM.N_508_cascade_\
        );

    \I__842\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5524\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__5524\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__839\ : CascadeMux
    port map (
            O => \N__5521\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__5518\,
            I => \U712_CHIP_RAM.N_477_cascade_\
        );

    \I__837\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5512\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5512\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\
        );

    \I__835\ : InMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__5506\,
            I => \U712_CHIP_RAM.N_406\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__5503\,
            I => \N__5500\
        );

    \I__832\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__830\ : Odrv4
    port map (
            O => \N__5494\,
            I => \U712_CHIP_RAM.N_430\
        );

    \I__829\ : InMux
    port map (
            O => \N__5491\,
            I => \N__5479\
        );

    \I__828\ : InMux
    port map (
            O => \N__5490\,
            I => \N__5479\
        );

    \I__827\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5479\
        );

    \I__826\ : InMux
    port map (
            O => \N__5488\,
            I => \N__5479\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5472\
        );

    \I__824\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5467\
        );

    \I__823\ : InMux
    port map (
            O => \N__5477\,
            I => \N__5467\
        );

    \I__822\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5462\
        );

    \I__821\ : InMux
    port map (
            O => \N__5475\,
            I => \N__5462\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__5472\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5467\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5462\,
            I => \U712_CHIP_RAM.N_44\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__816\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5449\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5449\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__814\ : CEMux
    port map (
            O => \N__5446\,
            I => \N__5442\
        );

    \I__813\ : CEMux
    port map (
            O => \N__5445\,
            I => \N__5439\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5436\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5433\
        );

    \I__810\ : Span4Mux_h
    port map (
            O => \N__5436\,
            I => \N__5430\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__5433\,
            I => \N__5427\
        );

    \I__808\ : Odrv4
    port map (
            O => \N__5430\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__5427\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__806\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5419\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5419\,
            I => \N__5415\
        );

    \I__804\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5412\
        );

    \I__803\ : Odrv4
    port map (
            O => \N__5415\,
            I => \U712_CHIP_RAM.N_500\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5412\,
            I => \U712_CHIP_RAM.N_500\
        );

    \I__801\ : InMux
    port map (
            O => \N__5407\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__800\ : InMux
    port map (
            O => \N__5404\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__799\ : InMux
    port map (
            O => \N__5401\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__798\ : InMux
    port map (
            O => \N__5398\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__797\ : ClkMux
    port map (
            O => \N__5395\,
            I => \N__5371\
        );

    \I__796\ : ClkMux
    port map (
            O => \N__5394\,
            I => \N__5371\
        );

    \I__795\ : ClkMux
    port map (
            O => \N__5393\,
            I => \N__5371\
        );

    \I__794\ : ClkMux
    port map (
            O => \N__5392\,
            I => \N__5371\
        );

    \I__793\ : ClkMux
    port map (
            O => \N__5391\,
            I => \N__5371\
        );

    \I__792\ : ClkMux
    port map (
            O => \N__5390\,
            I => \N__5371\
        );

    \I__791\ : ClkMux
    port map (
            O => \N__5389\,
            I => \N__5371\
        );

    \I__790\ : ClkMux
    port map (
            O => \N__5388\,
            I => \N__5371\
        );

    \I__789\ : GlobalMux
    port map (
            O => \N__5371\,
            I => \N__5368\
        );

    \I__788\ : gio2CtrlBuf
    port map (
            O => \N__5368\,
            I => \C1_c_g\
        );

    \I__787\ : SRMux
    port map (
            O => \N__5365\,
            I => \N__5362\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5362\,
            I => \N__5359\
        );

    \I__785\ : Odrv12
    port map (
            O => \N__5359\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__784\ : InMux
    port map (
            O => \N__5356\,
            I => \N__5352\
        );

    \I__783\ : InMux
    port map (
            O => \N__5355\,
            I => \N__5349\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5352\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5349\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__780\ : InMux
    port map (
            O => \N__5344\,
            I => \N__5340\
        );

    \I__779\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5337\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5340\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5337\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__776\ : InMux
    port map (
            O => \N__5332\,
            I => \N__5328\
        );

    \I__775\ : InMux
    port map (
            O => \N__5331\,
            I => \N__5325\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5328\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5325\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__772\ : InMux
    port map (
            O => \N__5320\,
            I => \N__5317\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__770\ : Odrv12
    port map (
            O => \N__5314\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\
        );

    \I__769\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__5305\,
            I => \N__5301\
        );

    \I__766\ : IoInMux
    port map (
            O => \N__5304\,
            I => \N__5298\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__5301\,
            I => \N__5295\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__5298\,
            I => \N__5292\
        );

    \I__763\ : Span4Mux_v
    port map (
            O => \N__5295\,
            I => \N__5289\
        );

    \I__762\ : IoSpan4Mux
    port map (
            O => \N__5292\,
            I => \N__5286\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__5289\,
            I => \RAMENn_c\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__5286\,
            I => \RAMENn_c\
        );

    \I__759\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5278\,
            I => \N__5274\
        );

    \I__757\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5271\
        );

    \I__756\ : Span4Mux_h
    port map (
            O => \N__5274\,
            I => \N__5266\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5271\,
            I => \N__5266\
        );

    \I__754\ : Span4Mux_v
    port map (
            O => \N__5266\,
            I => \N__5263\
        );

    \I__753\ : Sp12to4
    port map (
            O => \N__5263\,
            I => \N__5260\
        );

    \I__752\ : Span12Mux_h
    port map (
            O => \N__5260\,
            I => \N__5257\
        );

    \I__751\ : Odrv12
    port map (
            O => \N__5257\,
            I => \TSn_c\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__749\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__747\ : Odrv12
    port map (
            O => \N__5245\,
            I => \U712_CHIP_RAM.N_471\
        );

    \I__746\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5238\
        );

    \I__745\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5235\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5238\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5235\,
            I => \U712_CHIP_RAM.REFRESH5lto2\
        );

    \I__742\ : InMux
    port map (
            O => \N__5230\,
            I => \N__5226\
        );

    \I__741\ : InMux
    port map (
            O => \N__5229\,
            I => \N__5223\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__5226\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5223\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__738\ : CascadeMux
    port map (
            O => \N__5218\,
            I => \N__5214\
        );

    \I__737\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5211\
        );

    \I__736\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__5211\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5208\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__733\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5199\
        );

    \I__732\ : InMux
    port map (
            O => \N__5202\,
            I => \N__5196\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5199\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__5196\,
            I => \U712_CHIP_RAM.REFRESH5lto1\
        );

    \I__729\ : InMux
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__5185\,
            I => \N__5182\
        );

    \I__726\ : Odrv4
    port map (
            O => \N__5182\,
            I => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\
        );

    \I__725\ : IoInMux
    port map (
            O => \N__5179\,
            I => \N__5176\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5176\,
            I => \N__5173\
        );

    \I__723\ : Span4Mux_s2_v
    port map (
            O => \N__5173\,
            I => \N__5170\
        );

    \I__722\ : Span4Mux_v
    port map (
            O => \N__5170\,
            I => \N__5167\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__5167\,
            I => \N__5164\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__5164\,
            I => \VBENn_c\
        );

    \I__719\ : InMux
    port map (
            O => \N__5161\,
            I => \N__5158\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5158\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__717\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5151\
        );

    \I__716\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5143\
        );

    \I__714\ : InMux
    port map (
            O => \N__5150\,
            I => \N__5138\
        );

    \I__713\ : InMux
    port map (
            O => \N__5149\,
            I => \N__5138\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5146\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__5143\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5138\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__5131\,
            I => \U712_REG_SM.N_347_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__5125\,
            I => \U712_REG_SM.N_464\
        );

    \I__706\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__5119\,
            I => \U712_REG_SM.N_330\
        );

    \I__704\ : CascadeMux
    port map (
            O => \N__5116\,
            I => \U712_REG_SM.N_330_cascade_\
        );

    \I__703\ : InMux
    port map (
            O => \N__5113\,
            I => \bfn_9_15_0_\
        );

    \I__702\ : InMux
    port map (
            O => \N__5110\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__701\ : InMux
    port map (
            O => \N__5107\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__700\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5100\
        );

    \I__699\ : InMux
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5097\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__696\ : Odrv12
    port map (
            O => \N__5094\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__695\ : InMux
    port map (
            O => \N__5089\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5086\,
            I => \U712_CYCLE_TERM.N_486_cascade_\
        );

    \I__693\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5078\
        );

    \I__692\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5072\
        );

    \I__691\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5072\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5069\
        );

    \I__689\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5066\
        );

    \I__688\ : LocalMux
    port map (
            O => \N__5072\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__687\ : Odrv4
    port map (
            O => \N__5069\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5066\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__685\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5054\
        );

    \I__684\ : InMux
    port map (
            O => \N__5058\,
            I => \N__5049\
        );

    \I__683\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5049\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5054\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5049\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__679\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5038\,
            I => \U712_CYCLE_TERM.TACK_EN6_0\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__5035\,
            I => \U712_REG_SM.N_465_cascade_\
        );

    \I__676\ : InMux
    port map (
            O => \N__5032\,
            I => \N__5029\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5029\,
            I => \N__5026\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__5026\,
            I => \U712_CHIP_RAM.un3_DMA_CYCLE_START\
        );

    \I__673\ : CascadeMux
    port map (
            O => \N__5023\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__5020\,
            I => \U712_CHIP_RAM.N_402_cascade_\
        );

    \I__671\ : InMux
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__5014\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_3\
        );

    \I__669\ : InMux
    port map (
            O => \N__5011\,
            I => \N__5008\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__667\ : Span4Mux_v
    port map (
            O => \N__5005\,
            I => \N__5002\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__664\ : Sp12to4
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__4993\,
            I => \A_c_2\
        );

    \I__662\ : IoInMux
    port map (
            O => \N__4990\,
            I => \N__4987\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4987\,
            I => \N__4984\
        );

    \I__660\ : Span12Mux_s4_v
    port map (
            O => \N__4984\,
            I => \N__4980\
        );

    \I__659\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4977\
        );

    \I__658\ : Span12Mux_v
    port map (
            O => \N__4980\,
            I => \N__4972\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4977\,
            I => \N__4972\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__4972\,
            I => \N__4969\
        );

    \I__655\ : Odrv12
    port map (
            O => \N__4969\,
            I => \A_c_9\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__4966\,
            I => \U712_CHIP_RAM.REFRESH_RST_cascade_\
        );

    \I__653\ : CascadeMux
    port map (
            O => \N__4963\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__652\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4957\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4957\,
            I => \N__4954\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__4954\,
            I => \N__4951\
        );

    \I__649\ : Sp12to4
    port map (
            O => \N__4951\,
            I => \N__4948\
        );

    \I__648\ : Span12Mux_v
    port map (
            O => \N__4948\,
            I => \N__4945\
        );

    \I__647\ : Odrv12
    port map (
            O => \N__4945\,
            I => \A_c_14\
        );

    \I__646\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4939\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4939\,
            I => \N__4936\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__643\ : Sp12to4
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__642\ : Odrv12
    port map (
            O => \N__4930\,
            I => \A_c_7\
        );

    \I__641\ : CascadeMux
    port map (
            O => \N__4927\,
            I => \U712_CHIP_RAM.N_326_cascade_\
        );

    \I__640\ : InMux
    port map (
            O => \N__4924\,
            I => \N__4920\
        );

    \I__639\ : InMux
    port map (
            O => \N__4923\,
            I => \N__4917\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4914\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4909\
        );

    \I__636\ : Span4Mux_h
    port map (
            O => \N__4914\,
            I => \N__4909\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4909\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_a2_1\
        );

    \I__634\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4903\,
            I => \U712_CHIP_RAM.N_614\
        );

    \I__632\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4897\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\
        );

    \I__630\ : CascadeMux
    port map (
            O => \N__4894\,
            I => \U712_CHIP_RAM.N_614_cascade_\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__4891\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_3_1_cascade_\
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__4888\,
            I => \U712_CHIP_RAM.N_338_cascade_\
        );

    \I__627\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4881\
        );

    \I__626\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4878\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4881\,
            I => \N__4875\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4878\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__4875\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__4870\,
            I => \U712_CHIP_RAM.N_430_cascade_\
        );

    \I__621\ : InMux
    port map (
            O => \N__4867\,
            I => \N__4864\
        );

    \I__620\ : LocalMux
    port map (
            O => \N__4864\,
            I => \U712_CHIP_RAM.N_429\
        );

    \I__619\ : InMux
    port map (
            O => \N__4861\,
            I => \N__4856\
        );

    \I__618\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4851\
        );

    \I__617\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4851\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4856\,
            I => \N__4848\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4851\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__4848\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\
        );

    \I__613\ : InMux
    port map (
            O => \N__4843\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__612\ : InMux
    port map (
            O => \N__4840\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__611\ : InMux
    port map (
            O => \N__4837\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__610\ : InMux
    port map (
            O => \N__4834\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__609\ : InMux
    port map (
            O => \N__4831\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__608\ : InMux
    port map (
            O => \N__4828\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__607\ : InMux
    port map (
            O => \N__4825\,
            I => \N__4822\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4822\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_1\
        );

    \I__605\ : CascadeMux
    port map (
            O => \N__4819\,
            I => \U712_CHIP_RAM.N_515_cascade_\
        );

    \I__604\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4813\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__4813\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0\
        );

    \I__602\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4805\
        );

    \I__601\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4802\
        );

    \I__600\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4799\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4805\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4802\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4799\,
            I => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4792\,
            I => \U712_REG_SM.N_349_cascade_\
        );

    \I__595\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4786\,
            I => \U712_CHIP_RAM.CLK_EN_e_1\
        );

    \I__593\ : CascadeMux
    port map (
            O => \N__4783\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1_cascade_\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__4780\,
            I => \U712_CHIP_RAM.N_432_cascade_\
        );

    \I__591\ : InMux
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__4774\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \U712_CHIP_RAM.N_406_cascade_\
        );

    \I__588\ : InMux
    port map (
            O => \N__4768\,
            I => \bfn_9_7_0_\
        );

    \I__587\ : InMux
    port map (
            O => \N__4765\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__586\ : InMux
    port map (
            O => \N__4762\,
            I => \N__4758\
        );

    \I__585\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4755\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4758\,
            I => \N__4752\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__4755\,
            I => \N__4749\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4752\,
            I => \N__4746\
        );

    \I__581\ : Span4Mux_v
    port map (
            O => \N__4749\,
            I => \N__4743\
        );

    \I__580\ : Sp12to4
    port map (
            O => \N__4746\,
            I => \N__4740\
        );

    \I__579\ : Span4Mux_h
    port map (
            O => \N__4743\,
            I => \N__4737\
        );

    \I__578\ : Span12Mux_h
    port map (
            O => \N__4740\,
            I => \N__4732\
        );

    \I__577\ : Sp12to4
    port map (
            O => \N__4737\,
            I => \N__4732\
        );

    \I__576\ : Span12Mux_v
    port map (
            O => \N__4732\,
            I => \N__4729\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4729\,
            I => \DBRn_c\
        );

    \I__574\ : InMux
    port map (
            O => \N__4726\,
            I => \N__4723\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4723\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\
        );

    \I__572\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__571\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4714\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4714\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__569\ : IoInMux
    port map (
            O => \N__4711\,
            I => \N__4706\
        );

    \I__568\ : IoInMux
    port map (
            O => \N__4710\,
            I => \N__4703\
        );

    \I__567\ : IoInMux
    port map (
            O => \N__4709\,
            I => \N__4700\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4706\,
            I => \N__4697\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4703\,
            I => \N__4694\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4700\,
            I => \N__4691\
        );

    \I__563\ : Span4Mux_s3_v
    port map (
            O => \N__4697\,
            I => \N__4688\
        );

    \I__562\ : Span4Mux_s3_h
    port map (
            O => \N__4694\,
            I => \N__4685\
        );

    \I__561\ : Span12Mux_s4_v
    port map (
            O => \N__4691\,
            I => \N__4682\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__4688\,
            I => \N__4679\
        );

    \I__559\ : Span4Mux_h
    port map (
            O => \N__4685\,
            I => \N__4676\
        );

    \I__558\ : Span12Mux_h
    port map (
            O => \N__4682\,
            I => \N__4673\
        );

    \I__557\ : Span12Mux_s11_h
    port map (
            O => \N__4679\,
            I => \N__4670\
        );

    \I__556\ : Span4Mux_h
    port map (
            O => \N__4676\,
            I => \N__4667\
        );

    \I__555\ : Span12Mux_v
    port map (
            O => \N__4673\,
            I => \N__4663\
        );

    \I__554\ : Span12Mux_v
    port map (
            O => \N__4670\,
            I => \N__4658\
        );

    \I__553\ : Sp12to4
    port map (
            O => \N__4667\,
            I => \N__4658\
        );

    \I__552\ : InMux
    port map (
            O => \N__4666\,
            I => \N__4655\
        );

    \I__551\ : Odrv12
    port map (
            O => \N__4663\,
            I => \TACK_EN\
        );

    \I__550\ : Odrv12
    port map (
            O => \N__4658\,
            I => \TACK_EN\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4655\,
            I => \TACK_EN\
        );

    \I__548\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4643\
        );

    \I__547\ : InMux
    port map (
            O => \N__4647\,
            I => \N__4638\
        );

    \I__546\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4638\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__4643\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__4638\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__543\ : IoInMux
    port map (
            O => \N__4633\,
            I => \N__4630\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__4630\,
            I => \N__4626\
        );

    \I__541\ : IoInMux
    port map (
            O => \N__4629\,
            I => \N__4623\
        );

    \I__540\ : Span4Mux_s0_v
    port map (
            O => \N__4626\,
            I => \N__4619\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4623\,
            I => \N__4616\
        );

    \I__538\ : IoInMux
    port map (
            O => \N__4622\,
            I => \N__4613\
        );

    \I__537\ : Span4Mux_v
    port map (
            O => \N__4619\,
            I => \N__4610\
        );

    \I__536\ : IoSpan4Mux
    port map (
            O => \N__4616\,
            I => \N__4607\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4613\,
            I => \N__4604\
        );

    \I__534\ : Sp12to4
    port map (
            O => \N__4610\,
            I => \N__4601\
        );

    \I__533\ : Span4Mux_s2_v
    port map (
            O => \N__4607\,
            I => \N__4598\
        );

    \I__532\ : Span4Mux_s3_h
    port map (
            O => \N__4604\,
            I => \N__4595\
        );

    \I__531\ : Span12Mux_h
    port map (
            O => \N__4601\,
            I => \N__4592\
        );

    \I__530\ : Sp12to4
    port map (
            O => \N__4598\,
            I => \N__4589\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__4595\,
            I => \N__4586\
        );

    \I__528\ : Span12Mux_v
    port map (
            O => \N__4592\,
            I => \N__4578\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__4589\,
            I => \N__4578\
        );

    \I__526\ : Span12Mux_v
    port map (
            O => \N__4586\,
            I => \N__4578\
        );

    \I__525\ : InMux
    port map (
            O => \N__4585\,
            I => \N__4575\
        );

    \I__524\ : Odrv12
    port map (
            O => \N__4578\,
            I => \TACK_OUTn\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4575\,
            I => \TACK_OUTn\
        );

    \I__522\ : InMux
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4567\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__520\ : IoInMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__4561\,
            I => \N__4558\
        );

    \I__518\ : IoSpan4Mux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__517\ : Span4Mux_s1_v
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__516\ : Sp12to4
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__515\ : Span12Mux_v
    port map (
            O => \N__4549\,
            I => \N__4544\
        );

    \I__514\ : InMux
    port map (
            O => \N__4548\,
            I => \N__4541\
        );

    \I__513\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4538\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4544\,
            I => \REGENn_c\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4541\,
            I => \REGENn_c\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__4538\,
            I => \REGENn_c\
        );

    \I__509\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4528\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__4528\,
            I => \U712_REG_SM.REGENn_e_1\
        );

    \I__507\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4521\
        );

    \I__506\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4518\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4521\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__4518\,
            I => \U712_REG_SM.STATE_COUNTZ1Z_0\
        );

    \I__503\ : InMux
    port map (
            O => \N__4513\,
            I => \N__4509\
        );

    \I__502\ : InMux
    port map (
            O => \N__4512\,
            I => \N__4506\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4509\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4506\,
            I => \U712_REG_SM.START_RSTZ0\
        );

    \I__499\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4498\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4498\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__4495\,
            I => \U712_CHIP_RAM.N_480_cascade_\
        );

    \I__496\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4489\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__4489\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3\
        );

    \I__494\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4483\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4483\,
            I => \N__4480\
        );

    \I__492\ : Span12Mux_v
    port map (
            O => \N__4480\,
            I => \N__4477\
        );

    \I__491\ : Odrv12
    port map (
            O => \N__4477\,
            I => \A_c_5\
        );

    \I__490\ : InMux
    port map (
            O => \N__4474\,
            I => \N__4471\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__4471\,
            I => \N__4468\
        );

    \I__488\ : Span4Mux_v
    port map (
            O => \N__4468\,
            I => \N__4465\
        );

    \I__487\ : Span4Mux_h
    port map (
            O => \N__4465\,
            I => \N__4462\
        );

    \I__486\ : Span4Mux_h
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__4459\,
            I => \A_c_12\
        );

    \I__484\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4453\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4453\,
            I => \N__4450\
        );

    \I__482\ : Span4Mux_v
    port map (
            O => \N__4450\,
            I => \N__4447\
        );

    \I__481\ : Span4Mux_h
    port map (
            O => \N__4447\,
            I => \N__4444\
        );

    \I__480\ : Span4Mux_h
    port map (
            O => \N__4444\,
            I => \N__4441\
        );

    \I__479\ : Odrv4
    port map (
            O => \N__4441\,
            I => \A_c_8\
        );

    \I__478\ : InMux
    port map (
            O => \N__4438\,
            I => \N__4435\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4435\,
            I => \N__4432\
        );

    \I__476\ : Span12Mux_v
    port map (
            O => \N__4432\,
            I => \N__4429\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4429\,
            I => \A_c_15\
        );

    \I__474\ : IoInMux
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__4423\,
            I => \N__4420\
        );

    \I__472\ : IoSpan4Mux
    port map (
            O => \N__4420\,
            I => \N__4417\
        );

    \I__471\ : Span4Mux_s2_v
    port map (
            O => \N__4417\,
            I => \N__4414\
        );

    \I__470\ : Sp12to4
    port map (
            O => \N__4414\,
            I => \N__4411\
        );

    \I__469\ : Span12Mux_s8_v
    port map (
            O => \N__4411\,
            I => \N__4407\
        );

    \I__468\ : InMux
    port map (
            O => \N__4410\,
            I => \N__4404\
        );

    \I__467\ : Span12Mux_h
    port map (
            O => \N__4407\,
            I => \N__4399\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4404\,
            I => \N__4399\
        );

    \I__465\ : Span12Mux_v
    port map (
            O => \N__4399\,
            I => \N__4396\
        );

    \I__464\ : Odrv12
    port map (
            O => \N__4396\,
            I => \A_c_11\
        );

    \I__463\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4390\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__4390\,
            I => \N__4387\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__4387\,
            I => \N__4384\
        );

    \I__460\ : Span4Mux_v
    port map (
            O => \N__4384\,
            I => \N__4381\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__4381\,
            I => \N__4378\
        );

    \I__458\ : Span12Mux_h
    port map (
            O => \N__4378\,
            I => \N__4375\
        );

    \I__457\ : Odrv12
    port map (
            O => \N__4375\,
            I => \A_c_4\
        );

    \I__456\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__454\ : Span4Mux_v
    port map (
            O => \N__4366\,
            I => \N__4363\
        );

    \I__453\ : Sp12to4
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__452\ : Span12Mux_h
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__451\ : Span12Mux_v
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__450\ : Odrv12
    port map (
            O => \N__4354\,
            I => \A_c_16\
        );

    \I__449\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__447\ : Span12Mux_h
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__446\ : Span12Mux_v
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__445\ : Odrv12
    port map (
            O => \N__4339\,
            I => \A_c_18\
        );

    \I__444\ : CascadeMux
    port map (
            O => \N__4336\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\
        );

    \I__443\ : IoInMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__441\ : IoSpan4Mux
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__440\ : Span4Mux_s3_h
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__439\ : Span4Mux_v
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__438\ : Span4Mux_h
    port map (
            O => \N__4318\,
            I => \N__4315\
        );

    \I__437\ : Sp12to4
    port map (
            O => \N__4315\,
            I => \N__4311\
        );

    \I__436\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4308\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__4311\,
            I => \CLK_EN_c\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__4308\,
            I => \CLK_EN_c\
        );

    \I__433\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4300\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__4300\,
            I => \U712_CHIP_RAM.CLK_EN_6_0_a2_0_a2_1_0\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__4297\,
            I => \U712_CHIP_RAM.N_607_cascade_\
        );

    \I__430\ : InMux
    port map (
            O => \N__4294\,
            I => \N__4291\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4291\,
            I => \N__4288\
        );

    \I__428\ : Span4Mux_h
    port map (
            O => \N__4288\,
            I => \N__4285\
        );

    \I__427\ : Span4Mux_v
    port map (
            O => \N__4285\,
            I => \N__4282\
        );

    \I__426\ : Sp12to4
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4279\,
            I => \A_c_6\
        );

    \I__424\ : InMux
    port map (
            O => \N__4276\,
            I => \N__4273\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__422\ : Span12Mux_v
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__421\ : Odrv12
    port map (
            O => \N__4267\,
            I => \A_c_13\
        );

    \I__420\ : CascadeMux
    port map (
            O => \N__4264\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__418\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__4255\,
            I => \U712_CHIP_RAM.N_484\
        );

    \I__416\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4246\
        );

    \I__415\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4246\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4246\,
            I => \U712_CHIP_RAM.N_607\
        );

    \I__413\ : InMux
    port map (
            O => \N__4243\,
            I => \N__4237\
        );

    \I__412\ : InMux
    port map (
            O => \N__4242\,
            I => \N__4237\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4237\,
            I => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\
        );

    \I__410\ : InMux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4231\,
            I => \U712_REG_SM.N_456\
        );

    \I__408\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4224\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__4227\,
            I => \N__4221\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4224\,
            I => \N__4218\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4221\,
            I => \N__4215\
        );

    \I__404\ : Span4Mux_v
    port map (
            O => \N__4218\,
            I => \N__4212\
        );

    \I__403\ : IoSpan4Mux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__4212\,
            I => \N__4206\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__400\ : Span12Mux_h
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__399\ : IoSpan4Mux
    port map (
            O => \N__4203\,
            I => \N__4197\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__4200\,
            I => \C1_c\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__4197\,
            I => \C1_c\
        );

    \I__396\ : InMux
    port map (
            O => \N__4192\,
            I => \N__4189\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4189\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__394\ : InMux
    port map (
            O => \N__4186\,
            I => \N__4183\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__4183\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__392\ : IoInMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4177\,
            I => \N__4174\
        );

    \I__390\ : Span4Mux_s3_v
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__389\ : Span4Mux_v
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__388\ : Span4Mux_v
    port map (
            O => \N__4168\,
            I => \N__4164\
        );

    \I__387\ : InMux
    port map (
            O => \N__4167\,
            I => \N__4161\
        );

    \I__386\ : Odrv4
    port map (
            O => \N__4164\,
            I => \DBDIR_c\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__4161\,
            I => \DBDIR_c\
        );

    \I__384\ : IoInMux
    port map (
            O => \N__4156\,
            I => \N__4153\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__382\ : Odrv12
    port map (
            O => \N__4150\,
            I => \DBRn_c_i_0\
        );

    \I__381\ : IoInMux
    port map (
            O => \N__4147\,
            I => \N__4144\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__4144\,
            I => \N__4141\
        );

    \I__379\ : Span4Mux_s2_v
    port map (
            O => \N__4141\,
            I => \N__4138\
        );

    \I__378\ : Span4Mux_v
    port map (
            O => \N__4138\,
            I => \N__4135\
        );

    \I__377\ : Span4Mux_h
    port map (
            O => \N__4135\,
            I => \N__4132\
        );

    \I__376\ : Odrv4
    port map (
            O => \N__4132\,
            I => \CLK80_PLL_i_i\
        );

    \I__375\ : InMux
    port map (
            O => \N__4129\,
            I => \N__4126\
        );

    \I__374\ : LocalMux
    port map (
            O => \N__4126\,
            I => \N__4123\
        );

    \I__373\ : Span12Mux_h
    port map (
            O => \N__4123\,
            I => \N__4120\
        );

    \I__372\ : Span12Mux_v
    port map (
            O => \N__4120\,
            I => \N__4117\
        );

    \I__371\ : Odrv12
    port map (
            O => \N__4117\,
            I => \REGSPACEn_c\
        );

    \I__370\ : IoInMux
    port map (
            O => \N__4114\,
            I => \N__4111\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__4111\,
            I => \N__4108\
        );

    \I__368\ : IoSpan4Mux
    port map (
            O => \N__4108\,
            I => \N__4105\
        );

    \I__367\ : IoSpan4Mux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__366\ : Span4Mux_s3_h
    port map (
            O => \N__4102\,
            I => \N__4098\
        );

    \I__365\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4095\
        );

    \I__364\ : Span4Mux_h
    port map (
            O => \N__4098\,
            I => \N__4092\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__4095\,
            I => \N__4089\
        );

    \I__362\ : Sp12to4
    port map (
            O => \N__4092\,
            I => \N__4086\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__4089\,
            I => \N__4083\
        );

    \I__360\ : Span12Mux_h
    port map (
            O => \N__4086\,
            I => \N__4078\
        );

    \I__359\ : Sp12to4
    port map (
            O => \N__4083\,
            I => \N__4078\
        );

    \I__358\ : Span12Mux_h
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__357\ : Odrv12
    port map (
            O => \N__4075\,
            I => \C3_c\
        );

    \I__356\ : IoInMux
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__4069\,
            I => \N__4066\
        );

    \I__354\ : IoSpan4Mux
    port map (
            O => \N__4066\,
            I => \N__4063\
        );

    \I__353\ : Span4Mux_s2_v
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__352\ : Sp12to4
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__351\ : Span12Mux_v
    port map (
            O => \N__4057\,
            I => \N__4054\
        );

    \I__350\ : Odrv12
    port map (
            O => \N__4054\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            I => \N__5395\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            I => \N__5393\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__5394\
        );

    \INVU712_CHIP_RAM.DMA_A1_nesrC\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            I => \N__5390\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__5392\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__5388\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__5391\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_15_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4227\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__8647\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4156\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4114\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9267\,
            in2 => \_gnd_net_\,
            in3 => \N__10417\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9415\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4761\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5281\,
            in2 => \_gnd_net_\,
            in3 => \N__4129\,
            lcout => \U712_REG_SM.N_456\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4101\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9411\,
            ce => 'H',
            sr => \N__10368\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__9124\,
            in1 => \N__8838\,
            in2 => \_gnd_net_\,
            in3 => \N__5083\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4646\,
            in2 => \_gnd_net_\,
            in3 => \N__4242\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4243\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8839\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4647\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9401\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REGENn_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100011011000100"
        )
    port map (
            in0 => \N__4531\,
            in1 => \N__4548\,
            in2 => \N__9006\,
            in3 => \N__4525\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9404\,
            ce => 'H',
            sr => \N__10372\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__5150\,
            in1 => \N__4234\,
            in2 => \N__8857\,
            in3 => \N__4513\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9408\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5149\,
            in1 => \N__5897\,
            in2 => \N__8981\,
            in3 => \N__4524\,
            lcout => \U712_REG_SM.STATE_COUNT_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_0_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4228\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9410\,
            ce => 'H',
            sr => \N__10362\
        );

    \U712_REG_SM.C1_SYNC_1_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4192\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9410\,
            ce => 'H',
            sr => \N__10362\
        );

    \U712_REG_SM.C3_SYNC_1_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9410\,
            ce => 'H',
            sr => \N__10362\
        );

    \U712_REG_SM.WRITE_CYCLE_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__10261\,
            in1 => \N__5940\,
            in2 => \_gnd_net_\,
            in3 => \N__4808\,
            lcout => \U712_REG_SM.WRITE_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9410\,
            ce => 'H',
            sr => \N__10362\
        );

    \U712_CHIP_RAM.DBDIR_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4167\,
            in1 => \N__5722\,
            in2 => \_gnd_net_\,
            in3 => \N__6769\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => 'H',
            sr => \N__10394\
        );

    \U712_CHIP_RAM.CLK_EN_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__4789\,
            in1 => \N__4314\,
            in2 => \N__5611\,
            in3 => \N__4303\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9385\,
            ce => 'H',
            sr => \N__10394\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_0_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7271\,
            in1 => \N__6424\,
            in2 => \N__10200\,
            in3 => \N__7819\,
            lcout => \U712_CHIP_RAM.CLK_EN_6_0_a2_0_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR80N2_4_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6480\,
            lcout => \U712_CHIP_RAM.N_607\,
            ltout => \U712_CHIP_RAM.N_607_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__7270\,
            in1 => \N__6423\,
            in2 => \N__4297\,
            in3 => \N__7193\,
            lcout => \U712_CHIP_RAM.N_484\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4294\,
            in1 => \N__4276\,
            in2 => \_gnd_net_\,
            in3 => \N__8180\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIE24B8_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4924\,
            in1 => \N__4906\,
            in2 => \_gnd_net_\,
            in3 => \N__5596\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110000"
        )
    port map (
            in0 => \N__7328\,
            in1 => \N__7272\,
            in2 => \N__4264\,
            in3 => \N__4251\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001101"
        )
    port map (
            in0 => \N__4859\,
            in1 => \N__8181\,
            in2 => \N__4261\,
            in3 => \N__4816\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__4252\,
            in1 => \N__7329\,
            in2 => \N__7284\,
            in3 => \N__7198\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_480_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101100000001"
        )
    port map (
            in0 => \N__4860\,
            in1 => \N__4501\,
            in2 => \N__4495\,
            in3 => \N__6248\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9391\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__4861\,
            in1 => \N__4492\,
            in2 => \_gnd_net_\,
            in3 => \N__9878\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9393\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__8157\,
            in2 => \_gnd_net_\,
            in3 => \N__4474\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4456\,
            in1 => \N__4438\,
            in2 => \_gnd_net_\,
            in3 => \N__8156\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6611\,
            in1 => \N__9618\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4410\,
            in1 => \N__4393\,
            in2 => \_gnd_net_\,
            in3 => \N__8155\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIHJRU1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__8814\,
            in1 => \N__6600\,
            in2 => \N__9617\,
            in3 => \N__6569\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4372\,
            in1 => \N__4351\,
            in2 => \_gnd_net_\,
            in3 => \N__8189\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8190\,
            in1 => \N__7818\,
            in2 => \N__4336\,
            in3 => \N__10795\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4762\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => 'H',
            sr => \N__10373\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__4726\,
            in1 => \N__4720\,
            in2 => \N__5044\,
            in3 => \N__5081\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => 'H',
            sr => \N__10373\
        );

    \U712_CYCLE_TERM.TACK_EN_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011111111"
        )
    port map (
            in0 => \N__4719\,
            in1 => \N__4666\,
            in2 => \_gnd_net_\,
            in3 => \N__5632\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => 'H',
            sr => \N__10373\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110110011101110"
        )
    port map (
            in0 => \N__4585\,
            in1 => \N__4648\,
            in2 => \N__9131\,
            in3 => \N__5082\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => 'H',
            sr => \N__10373\
        );

    \DBR_SYNC_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4570\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9398\,
            ce => 'H',
            sr => \N__10373\
        );

    \U712_REG_SM.REGENn_RNO_0_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001011000"
        )
    port map (
            in0 => \N__4547\,
            in1 => \N__6017\,
            in2 => \N__5919\,
            in3 => \N__5154\,
            lcout => \U712_REG_SM.REGENn_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_0_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__6058\,
            in1 => \N__5122\,
            in2 => \N__5848\,
            in3 => \N__5128\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__10363\
        );

    \U712_REG_SM.START_RST_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__4512\,
            in1 => \N__4809\,
            in2 => \_gnd_net_\,
            in3 => \N__6009\,
            lcout => \U712_REG_SM.START_RSTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9405\,
            ce => 'H',
            sr => \N__10363\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5901\,
            in2 => \_gnd_net_\,
            in3 => \N__8959\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_349_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__8813\,
            in1 => \N__4810\,
            in2 => \N__4792\,
            in3 => \N__6010\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9409\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_RNO_1_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6454\,
            in1 => \N__6849\,
            in2 => \N__7192\,
            in3 => \N__6737\,
            lcout => \U712_CHIP_RAM.CLK_EN_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_3_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__7169\,
            in1 => \_gnd_net_\,
            in2 => \N__7278\,
            in3 => \N__7304\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIU95J5_4_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101000000000"
        )
    port map (
            in0 => \N__9746\,
            in1 => \N__6535\,
            in2 => \N__4783\,
            in3 => \N__9545\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITIV55_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__6453\,
            in1 => \N__5763\,
            in2 => \N__7191\,
            in3 => \N__6736\,
            lcout => \U712_CHIP_RAM.N_432\,
            ltout => \U712_CHIP_RAM.N_432_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJSRL5_0_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__8844\,
            in1 => \_gnd_net_\,
            in2 => \N__4780\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_406\,
            ltout => \U712_CHIP_RAM.N_406_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIHBUSE_4_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__4777\,
            in1 => \N__5422\,
            in2 => \N__4771\,
            in3 => \N__6484\,
            lcout => \U712_CHIP_RAM.N_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7178\,
            in2 => \_gnd_net_\,
            in3 => \N__4768\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5488\,
            in1 => \N__6848\,
            in2 => \_gnd_net_\,
            in3 => \N__4765\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6405\,
            in2 => \_gnd_net_\,
            in3 => \N__4843\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5489\,
            in1 => \N__7276\,
            in2 => \_gnd_net_\,
            in3 => \N__4840\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5475\,
            in1 => \N__6536\,
            in2 => \_gnd_net_\,
            in3 => \N__4837\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5490\,
            in1 => \N__5551\,
            in2 => \_gnd_net_\,
            in3 => \N__4834\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5476\,
            in1 => \N__5563\,
            in2 => \_gnd_net_\,
            in3 => \N__4831\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__5491\,
            in1 => \N__5575\,
            in2 => \_gnd_net_\,
            in3 => \N__4828\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9386\,
            ce => \N__5446\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_4_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__9534\,
            in1 => \_gnd_net_\,
            in2 => \N__6539\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_515\,
            ltout => \U712_CHIP_RAM.N_515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__4825\,
            in1 => \N__5801\,
            in2 => \N__4819\,
            in3 => \N__4923\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_58_i_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_2_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000110000"
        )
    port map (
            in0 => \N__7258\,
            in1 => \N__6398\,
            in2 => \N__6855\,
            in3 => \N__7156\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_326_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIBOVM2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__9690\,
            in1 => \_gnd_net_\,
            in2 => \N__4927\,
            in3 => \N__8817\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_134_i_a2_0_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6538\,
            in3 => \N__9689\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERlde_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_2_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9756\,
            in1 => \N__9535\,
            in2 => \_gnd_net_\,
            in3 => \N__8819\,
            lcout => \U712_CHIP_RAM.N_614\,
            ltout => \U712_CHIP_RAM.N_614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4TF5A_4_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__5802\,
            in1 => \N__4900\,
            in2 => \N__4894\,
            in3 => \N__4885\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIMEP34_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__7157\,
            in1 => \N__8818\,
            in2 => \N__6865\,
            in3 => \N__6727\,
            lcout => \U712_CHIP_RAM.N_429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_3_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__7185\,
            in1 => \N__6861\,
            in2 => \_gnd_net_\,
            in3 => \N__7279\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_a2_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIQGOH4_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__5418\,
            in1 => \N__9694\,
            in2 => \N__4891\,
            in3 => \N__9536\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIGCGV5_4_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6541\,
            in1 => \N__8815\,
            in2 => \N__4888\,
            in3 => \N__6416\,
            lcout => \U712_CHIP_RAM.N_430\,
            ltout => \U712_CHIP_RAM.N_430_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNILH2MF_1_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__4884\,
            in1 => \N__5800\,
            in2 => \N__4870\,
            in3 => \N__4867\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__5017\,
            in1 => \N__5740\,
            in2 => \N__5023\,
            in3 => \N__9826\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9392\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__7280\,
            in1 => \N__9695\,
            in2 => \N__7330\,
            in3 => \N__7186\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_402_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__9696\,
            in1 => \N__5734\,
            in2 => \N__5020\,
            in3 => \N__6417\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIR9VE1_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6601\,
            in1 => \N__5058\,
            in2 => \N__6096\,
            in3 => \N__9599\,
            lcout => \U712_CHIP_RAM.N_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__8188\,
            in1 => \N__5011\,
            in2 => \_gnd_net_\,
            in3 => \N__4983\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__6249\,
            in1 => \N__9871\,
            in2 => \N__9827\,
            in3 => \N__8185\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => \U712_CHIP_RAM.REFRESH_RST_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__8186\,
            in1 => \N__9872\,
            in2 => \N__4966\,
            in3 => \N__6250\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10416\,
            in1 => \_gnd_net_\,
            in2 => \N__4963\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8187\,
            in1 => \N__4960\,
            in2 => \_gnd_net_\,
            in3 => \N__4942\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5057\,
            in2 => \_gnd_net_\,
            in3 => \N__6083\,
            lcout => \U712_CHIP_RAM.N_327\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100110011"
        )
    port map (
            in0 => \N__6045\,
            in1 => \N__5077\,
            in2 => \N__5680\,
            in3 => \N__5649\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__5650\,
            in1 => \N__9132\,
            in2 => \N__5086\,
            in3 => \N__8699\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010110000"
        )
    port map (
            in0 => \N__5104\,
            in1 => \N__5320\,
            in2 => \N__8743\,
            in3 => \N__5191\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110001000"
        )
    port map (
            in0 => \N__8695\,
            in1 => \N__5032\,
            in2 => \N__9475\,
            in3 => \N__9610\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001010100000"
        )
    port map (
            in0 => \N__8694\,
            in1 => \N__7811\,
            in2 => \N__5254\,
            in3 => \N__5059\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9394\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6044\,
            in2 => \_gnd_net_\,
            in3 => \N__5676\,
            lcout => \U712_CYCLE_TERM.TACK_EN6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__5841\,
            in1 => \N__6950\,
            in2 => \_gnd_net_\,
            in3 => \N__6927\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_465_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__8810\,
            in1 => \N__5920\,
            in2 => \N__5035\,
            in3 => \N__9005\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9399\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5161\,
            in2 => \_gnd_net_\,
            in3 => \N__6906\,
            lcout => \U712_CHIP_RAM.un3_DMA_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6907\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8811\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9402\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNINRSB_2_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6949\,
            in2 => \_gnd_net_\,
            in3 => \N__6008\,
            lcout => \U712_REG_SM.N_347\,
            ltout => \U712_REG_SM.N_347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5155\,
            in1 => \N__5840\,
            in2 => \N__5131\,
            in3 => \N__5969\,
            lcout => \U712_REG_SM.N_464\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_0_4_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011101110"
        )
    port map (
            in0 => \N__5967\,
            in1 => \N__5910\,
            in2 => \_gnd_net_\,
            in3 => \N__8970\,
            lcout => \U712_REG_SM.N_330\,
            ltout => \U712_REG_SM.N_330_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_4_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__5847\,
            in1 => \N__8812\,
            in2 => \N__5116\,
            in3 => \N__5968\,
            lcout => \U712_REG_SM.STATE_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9406\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5230\,
            in2 => \_gnd_net_\,
            in3 => \N__5113\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_9_15_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5203\,
            in2 => \_gnd_net_\,
            in3 => \N__5110\,
            lcout => \U712_CHIP_RAM.REFRESH5lto1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5242\,
            in2 => \_gnd_net_\,
            in3 => \N__5107\,
            lcout => \U712_CHIP_RAM.REFRESH5lto2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5103\,
            in2 => \_gnd_net_\,
            in3 => \N__5089\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5217\,
            in2 => \_gnd_net_\,
            in3 => \N__5407\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5332\,
            in2 => \_gnd_net_\,
            in3 => \N__5404\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5344\,
            in2 => \_gnd_net_\,
            in3 => \N__5401\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5356\,
            in2 => \_gnd_net_\,
            in3 => \N__5398\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5389\,
            ce => 'H',
            sr => \N__5365\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5355\,
            in1 => \N__5343\,
            in2 => \_gnd_net_\,
            in3 => \N__5331\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5311\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5277\,
            lcout => \U712_CHIP_RAM.N_471\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111101011111"
        )
    port map (
            in0 => \N__5241\,
            in1 => \N__5229\,
            in2 => \N__5218\,
            in3 => \N__5202\,
            lcout => \U712_CHIP_RAM.REFRESH_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_0_a2_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7817\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11067\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_2_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6391\,
            in2 => \_gnd_net_\,
            in3 => \N__6851\,
            lcout => \U712_CHIP_RAM.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_1_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7809\,
            in1 => \N__7087\,
            in2 => \N__10195\,
            in3 => \N__5604\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__6852\,
            in1 => \N__7810\,
            in2 => \N__5518\,
            in3 => \N__10185\,
            lcout => \CPU_TACKm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9380\,
            ce => \N__6883\,
            sr => \N__10390\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIQTMR1_0_2_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6850\,
            in1 => \N__7252\,
            in2 => \N__6406\,
            in3 => \N__7152\,
            lcout => \U712_CHIP_RAM.N_501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001110101010"
        )
    port map (
            in0 => \N__5515\,
            in1 => \N__5509\,
            in2 => \N__5503\,
            in3 => \N__5478\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9382\,
            ce => \N__5445\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_RNO_0_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9748\,
            in1 => \N__9538\,
            in2 => \_gnd_net_\,
            in3 => \N__10951\,
            lcout => \U712_CHIP_RAM.DBENn_8_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIURFN4_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9537\,
            in1 => \N__9747\,
            in2 => \_gnd_net_\,
            in3 => \N__5782\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__5477\,
            in1 => \N__8855\,
            in2 => \N__5455\,
            in3 => \N__5530\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9382\,
            ce => \N__5445\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIR5PC1_0_3_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7155\,
            in1 => \N__6832\,
            in2 => \_gnd_net_\,
            in3 => \N__7254\,
            lcout => \U712_CHIP_RAM.N_500\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011100000"
        )
    port map (
            in0 => \N__10162\,
            in1 => \N__6392\,
            in2 => \N__6854\,
            in3 => \N__7153\,
            lcout => \U712_CHIP_RAM.N_608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__8837\,
            in1 => \N__9692\,
            in2 => \N__5623\,
            in3 => \N__5603\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9387\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5574\,
            in1 => \N__5562\,
            in2 => \_gnd_net_\,
            in3 => \N__5550\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5O1M2_4_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__6522\,
            in1 => \N__7253\,
            in2 => \N__5539\,
            in3 => \N__9691\,
            lcout => \U712_CHIP_RAM.N_504\,
            ltout => \U712_CHIP_RAM.N_504_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIN38L4_2_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6397\,
            in2 => \N__5536\,
            in3 => \N__5756\,
            lcout => \U712_CHIP_RAM.N_438\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIJJ8G1_0_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__7154\,
            in1 => \N__10163\,
            in2 => \N__6407\,
            in3 => \N__6831\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8HNG_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6393\,
            in2 => \_gnd_net_\,
            in3 => \N__9450\,
            lcout => \U712_CHIP_RAM.N_341\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIU2TJ3_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9755\,
            in1 => \N__9687\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \U712_CHIP_RAM.N_508\,
            ltout => \U712_CHIP_RAM.N_508_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIPCS25_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010110000"
        )
    port map (
            in0 => \N__9619\,
            in1 => \N__6619\,
            in2 => \N__5533\,
            in3 => \N__6570\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__8836\,
            in1 => \N__10173\,
            in2 => \N__5521\,
            in3 => \N__5686\,
            lcout => \WRITE_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNO_0_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5803\,
            in1 => \N__5781\,
            in2 => \N__5767\,
            in3 => \N__6735\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000001000"
        )
    port map (
            in0 => \N__8834\,
            in1 => \N__7776\,
            in2 => \N__5743\,
            in3 => \N__6121\,
            lcout => \CPU_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9389\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101001111"
        )
    port map (
            in0 => \N__10167\,
            in1 => \N__9688\,
            in2 => \N__9550\,
            in3 => \N__7190\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_3_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100110011"
        )
    port map (
            in0 => \N__6540\,
            in1 => \N__8835\,
            in2 => \_gnd_net_\,
            in3 => \N__6853\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_28_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__5728\,
            in1 => \N__7761\,
            in2 => \N__8257\,
            in3 => \N__10711\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6260\,
            in2 => \_gnd_net_\,
            in3 => \N__9820\,
            lcout => \U712_CHIP_RAM.N_337\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__9606\,
            in1 => \N__10269\,
            in2 => \_gnd_net_\,
            in3 => \N__5721\,
            lcout => \U712_CHIP_RAM.N_361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__6043\,
            in1 => \N__5675\,
            in2 => \_gnd_net_\,
            in3 => \N__5648\,
            lcout => \U712_CYCLE_TERM.N_350\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111011"
        )
    port map (
            in0 => \N__5918\,
            in1 => \N__6019\,
            in2 => \N__9007\,
            in3 => \N__6951\,
            lcout => \U712_REG_SM.STATE_COUNTc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5917\,
            in2 => \_gnd_net_\,
            in3 => \N__6097\,
            lcout => \U712_REG_SM.N_348\,
            ltout => \U712_REG_SM.N_348_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_2_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100000000"
        )
    port map (
            in0 => \N__8994\,
            in1 => \N__6067\,
            in2 => \N__6061\,
            in3 => \N__8833\,
            lcout => \U712_REG_SM.STATE_COUNTZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9395\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CUUBEn_i_0_a2_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011100000000"
        )
    port map (
            in0 => \N__7657\,
            in1 => \N__8520\,
            in2 => \N__8356\,
            in3 => \N__7816\,
            lcout => \U712_BYTE_ENABLE.N_441\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__6057\,
            in1 => \N__5809\,
            in2 => \N__6046\,
            in3 => \N__5926\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9400\,
            ce => 'H',
            sr => \N__10359\
        );

    \U712_REG_SM.STATE_COUNT_RNIVCF31_4_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100111"
        )
    port map (
            in0 => \N__8963\,
            in1 => \N__5970\,
            in2 => \N__6018\,
            in3 => \N__5902\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNT_RNIKVGT_4_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__5971\,
            in1 => \N__5908\,
            in2 => \_gnd_net_\,
            in3 => \N__8964\,
            lcout => \U712_REG_SM.N_399\,
            ltout => \U712_REG_SM.N_399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__5846\,
            in1 => \_gnd_net_\,
            in2 => \N__5944\,
            in3 => \N__5941\,
            lcout => \U712_REG_SM.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__8971\,
            in1 => \N__5909\,
            in2 => \_gnd_net_\,
            in3 => \N__5845\,
            lcout => \U712_REG_SM.N_458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011111010"
        )
    port map (
            in0 => \N__6325\,
            in1 => \N__6336\,
            in2 => \N__9008\,
            in3 => \N__7428\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9407\,
            ce => 'H',
            sr => \N__10355\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000100000"
        )
    port map (
            in0 => \N__8483\,
            in1 => \N__10262\,
            in2 => \N__8588\,
            in3 => \N__8398\,
            lcout => \U712_REG_SM.N_447\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.RASn_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6265\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9372\,
            ce => 'H',
            sr => \N__10391\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__6307\,
            in2 => \N__7831\,
            in3 => \N__10492\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9378\,
            ce => \N__7930\,
            sr => \N__10388\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__6261\,
            in1 => \N__8238\,
            in2 => \_gnd_net_\,
            in3 => \N__9834\,
            lcout => \U712_CHIP_RAM.CMA_5_i_0_8\,
            ltout => \U712_CHIP_RAM.CMA_5_i_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__6211\,
            in1 => \N__7812\,
            in2 => \N__6190\,
            in3 => \N__9772\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9378\,
            ce => \N__7930\,
            sr => \N__10388\
        );

    \U712_CHIP_RAM.BANK0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001011111110"
        )
    port map (
            in0 => \N__6132\,
            in1 => \N__6547\,
            in2 => \N__6163\,
            in3 => \N__6103\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9381\,
            ce => 'H',
            sr => \N__10383\
        );

    \U712_CHIP_RAM.BANK0_RNO_4_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9638\,
            in1 => \N__9750\,
            in2 => \_gnd_net_\,
            in3 => \N__9528\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.BANK0_RNOZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_1_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__6961\,
            in1 => \N__6117\,
            in2 => \N__6106\,
            in3 => \N__9253\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_2_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000000"
        )
    port map (
            in0 => \N__6618\,
            in1 => \N__6574\,
            in2 => \N__9640\,
            in3 => \N__9749\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_8_0_0_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6550\,
            in3 => \N__6479\,
            lcout => \U712_CHIP_RAM.N_433\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI5V372_4_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6537\,
            in1 => \N__9686\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \U712_CHIP_RAM.N_499\,
            ltout => \U712_CHIP_RAM.N_499_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_4_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7303\,
            in2 => \N__6457\,
            in3 => \N__7277\,
            lcout => \U712_CHIP_RAM.N_439\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6726\,
            in1 => \N__7177\,
            in2 => \N__6871\,
            in3 => \N__6452\,
            lcout => \U712_CHIP_RAM.N_507\,
            ltout => \U712_CHIP_RAM.N_507_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIALFTC_2_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6761\,
            in2 => \N__6436\,
            in3 => \N__6433\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__10415\,
            in1 => \_gnd_net_\,
            in2 => \N__6427\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9754\,
            in1 => \N__9693\,
            in2 => \N__9634\,
            in3 => \N__9529\,
            lcout => \U712_CHIP_RAM.BANK0_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_5_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6404\,
            in1 => \N__7176\,
            in2 => \N__6738\,
            in3 => \N__6869\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_440_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_2_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__6688\,
            in1 => \N__6731\,
            in2 => \N__6895\,
            in3 => \N__6892\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6886\,
            in3 => \N__10414\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6870\,
            in2 => \_gnd_net_\,
            in3 => \N__9470\,
            lcout => \U712_CHIP_RAM.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_RNO_1_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__6762\,
            in1 => \N__6745\,
            in2 => \N__6739\,
            in3 => \N__6687\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER46_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_CLK_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100010101000"
        )
    port map (
            in0 => \N__8845\,
            in1 => \N__6645\,
            in2 => \N__6673\,
            in3 => \N__6670\,
            lcout => \LATCH_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9388\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_RNI8NM9_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8227\,
            in2 => \_gnd_net_\,
            in3 => \N__7756\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_RNI8NMZ0Z9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110001111"
        )
    port map (
            in0 => \N__7980\,
            in1 => \N__9228\,
            in2 => \N__8253\,
            in3 => \N__7757\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000110011"
        )
    port map (
            in0 => \N__9229\,
            in1 => \N__8236\,
            in2 => \N__7808\,
            in3 => \N__7981\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6634\,
            in2 => \N__6628\,
            in3 => \N__6625\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9390\,
            ce => \N__7915\,
            sr => \N__10364\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8042\,
            in1 => \N__9967\,
            in2 => \N__7997\,
            in3 => \N__7039\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9390\,
            ce => \N__7915\,
            sr => \N__10364\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a2_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011110000"
        )
    port map (
            in0 => \N__8355\,
            in1 => \N__9028\,
            in2 => \N__7832\,
            in3 => \N__7654\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_443_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_32_i_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9195\,
            in1 => \N__10114\,
            in2 => \N__7009\,
            in3 => \N__9474\,
            lcout => \N_32_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_RNO_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10698\,
            in2 => \_gnd_net_\,
            in3 => \N__6982\,
            lcout => \U712_CHIP_RAM.BANK0_RNOZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6952\,
            in1 => \N__6928\,
            in2 => \_gnd_net_\,
            in3 => \N__8995\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_462_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__8832\,
            in1 => \N__11054\,
            in2 => \N__6916\,
            in3 => \N__6913\,
            lcout => \REG_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__8823\,
            in1 => \N__10113\,
            in2 => \_gnd_net_\,
            in3 => \N__11134\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9396\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_x2_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__8590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8443\,
            lcout => \U712_BYTE_ENABLE.N_323_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_RNO_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10413\,
            in2 => \_gnd_net_\,
            in3 => \N__7427\,
            lcout => \U712_REG_SM.un1_REGENn_0_sqmuxa_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1011101110111000"
        )
    port map (
            in0 => \N__7395\,
            in1 => \N__7429\,
            in2 => \N__9009\,
            in3 => \N__7384\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9403\,
            ce => 'H',
            sr => \N__10354\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10260\,
            in1 => \N__8484\,
            in2 => \N__8589\,
            in3 => \N__8445\,
            lcout => \U712_REG_SM.N_446\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DMA_LATCH_EN_i_i_a2_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__11123\,
            in1 => \N__10101\,
            in2 => \_gnd_net_\,
            in3 => \N__10196\,
            lcout => \N_435\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8254\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9370\,
            ce => 'H',
            sr => \N__10389\
        );

    \U712_CHIP_RAM.CPU_TACK_esr_RNO_3_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7311\,
            in1 => \N__7285\,
            in2 => \_gnd_net_\,
            in3 => \N__7197\,
            lcout => \U712_CHIP_RAM.CPU_TACK_7_iv_i_0_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DBENn_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__9172\,
            in1 => \N__7078\,
            in2 => \_gnd_net_\,
            in3 => \N__7072\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9374\,
            ce => 'H',
            sr => \N__10371\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__7820\,
            in1 => \N__7063\,
            in2 => \N__8255\,
            in3 => \N__10048\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__8014\,
            in1 => \N__8046\,
            in2 => \N__7627\,
            in3 => \N__10036\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9379\,
            ce => \N__7926\,
            sr => \N__10367\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000101"
        )
    port map (
            in0 => \N__8013\,
            in1 => \N__7477\,
            in2 => \N__8256\,
            in3 => \N__7450\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9379\,
            ce => \N__7926\,
            sr => \N__10367\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__8245\,
            in1 => \N__8016\,
            in2 => \_gnd_net_\,
            in3 => \N__9892\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9379\,
            ce => \N__7926\,
            sr => \N__10367\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100001000000"
        )
    port map (
            in0 => \N__8047\,
            in1 => \N__8015\,
            in2 => \N__7537\,
            in3 => \N__9217\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9379\,
            ce => \N__7926\,
            sr => \N__10367\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000010000"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__8237\,
            in2 => \N__10849\,
            in3 => \N__7546\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__8228\,
            in1 => \N__7806\,
            in2 => \N__7528\,
            in3 => \N__9985\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7803\,
            in1 => \N__7506\,
            in2 => \_gnd_net_\,
            in3 => \N__9916\,
            lcout => \U712_CHIP_RAM.N_382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__7471\,
            in1 => \N__7807\,
            in2 => \_gnd_net_\,
            in3 => \N__9976\,
            lcout => \U712_CHIP_RAM.N_374\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__7805\,
            in1 => \N__8229\,
            in2 => \N__7444\,
            in3 => \N__10858\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8266\,
            in1 => \N__7821\,
            in2 => \N__8252\,
            in3 => \N__10054\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010100000100000"
        )
    port map (
            in0 => \N__8008\,
            in1 => \N__8043\,
            in2 => \N__8098\,
            in3 => \N__9235\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__7925\,
            sr => \N__10360\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__8045\,
            in1 => \N__9958\,
            in2 => \N__8017\,
            in3 => \N__8071\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__7925\,
            sr => \N__10360\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010010000000"
        )
    port map (
            in0 => \N__8044\,
            in1 => \N__8012\,
            in2 => \N__9904\,
            in3 => \N__7960\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9384\,
            ce => \N__7925\,
            sr => \N__10360\
        );

    \U712_BYTE_ENABLE.N_34_i_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__9188\,
            in1 => \N__11133\,
            in2 => \N__7897\,
            in3 => \N__9473\,
            lcout => \N_34_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011110000"
        )
    port map (
            in0 => \N__8343\,
            in1 => \N__8524\,
            in2 => \N__7834\,
            in3 => \N__7656\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_451_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_200_i_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__9186\,
            in1 => \N__11132\,
            in2 => \N__7861\,
            in3 => \N__9471\,
            lcout => \N_200_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011110000"
        )
    port map (
            in0 => \N__8342\,
            in1 => \N__9027\,
            in2 => \N__7833\,
            in3 => \N__7655\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_453_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_202_i_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000001111"
        )
    port map (
            in0 => \N__9187\,
            in1 => \N__10089\,
            in2 => \N__9157\,
            in3 => \N__9472\,
            lcout => \N_202_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_RNI8MQ3_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_6_i_o2_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8449\,
            in2 => \_gnd_net_\,
            in3 => \N__8519\,
            lcout => \N_334\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.ASn_ess_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9010\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9397\,
            ce => \N__8872\,
            sr => \N__10353\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8786\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_353_i_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100110000"
        )
    port map (
            in0 => \N__8509\,
            in1 => \N__8314\,
            in2 => \N__8444\,
            in3 => \N__8569\,
            lcout => \N_353_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_354_i_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011000100"
        )
    port map (
            in0 => \N__8510\,
            in1 => \N__8566\,
            in2 => \N__8344\,
            in3 => \N__8417\,
            lcout => \N_354_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_84_i_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__8512\,
            in1 => \N__8568\,
            in2 => \N__8345\,
            in3 => \N__8421\,
            lcout => \N_84_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_355_i_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100001011010"
        )
    port map (
            in0 => \N__8567\,
            in1 => \N__8511\,
            in2 => \N__8433\,
            in3 => \N__8333\,
            lcout => \N_355_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CRCSn_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9891\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9371\,
            ce => 'H',
            sr => \N__10395\
        );

    \U712_CHIP_RAM.WEn_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9838\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9373\,
            ce => 'H',
            sr => \N__10392\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10834\,
            in1 => \N__10546\,
            in2 => \_gnd_net_\,
            in3 => \N__10693\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10477\,
            ce => \N__10452\,
            sr => \N__10384\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9760\,
            in1 => \N__9700\,
            in2 => \N__9639\,
            in3 => \N__9549\,
            lcout => \DMA_CYCLEm\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9383\,
            ce => \N__9286\,
            sr => \N__10374\
        );

    \U712_CHIP_RAM.DMA_A20_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__9274\,
            in1 => \N__10545\,
            in2 => \N__10699\,
            in3 => \N__9249\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10369\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__11023\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10475\,
            ce => \N__10448\,
            sr => \N__10365\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10782\,
            in1 => \N__10027\,
            in2 => \_gnd_net_\,
            in3 => \N__10666\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10475\,
            ce => \N__10448\,
            sr => \N__10365\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10667\,
            in1 => \N__10783\,
            in2 => \_gnd_net_\,
            in3 => \N__10747\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10475\,
            ce => \N__10448\,
            sr => \N__10365\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10673\,
            in1 => \N__11018\,
            in2 => \_gnd_net_\,
            in3 => \N__9947\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10446\,
            sr => \N__10361\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__10781\,
            in1 => \N__10674\,
            in2 => \_gnd_net_\,
            in3 => \N__10023\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__10446\,
            sr => \N__10361\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10022\,
            in1 => \N__10939\,
            in2 => \_gnd_net_\,
            in3 => \N__10689\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10476\,
            ce => \N__10453\,
            sr => \N__10385\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10021\,
            in1 => \N__10938\,
            in2 => \_gnd_net_\,
            in3 => \N__10688\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10450\,
            sr => \N__10375\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10687\,
            in1 => \N__9946\,
            in2 => \_gnd_net_\,
            in3 => \N__10892\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__10450\,
            sr => \N__10375\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10833\,
            in1 => \N__10746\,
            in2 => \_gnd_net_\,
            in3 => \N__10686\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10474\,
            ce => \N__10449\,
            sr => \N__10370\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9949\,
            in1 => \_gnd_net_\,
            in2 => \N__10697\,
            in3 => \N__10893\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10474\,
            ce => \N__10449\,
            sr => \N__10370\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__11019\,
            in1 => \N__9948\,
            in2 => \_gnd_net_\,
            in3 => \N__10681\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10474\,
            ce => \N__10449\,
            sr => \N__10370\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10894\,
            in1 => \N__10937\,
            in2 => \_gnd_net_\,
            in3 => \N__10685\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10474\,
            ce => \N__10449\,
            sr => \N__10370\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__11008\,
            in1 => \N__10980\,
            in2 => \_gnd_net_\,
            in3 => \N__10598\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A1_nesrC_net\,
            ce => \N__10447\,
            sr => \N__10366\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10927\,
            in1 => \N__10886\,
            in2 => \_gnd_net_\,
            in3 => \N__10680\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__10454\,
            sr => \N__10386\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10831\,
            in1 => \N__10745\,
            in2 => \_gnd_net_\,
            in3 => \N__10678\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10451\,
            sr => \N__10376\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10679\,
            in1 => \N__10832\,
            in2 => \_gnd_net_\,
            in3 => \N__10537\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6C_net\,
            ce => \N__10451\,
            sr => \N__10376\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10772\,
            in1 => \N__10744\,
            in2 => \_gnd_net_\,
            in3 => \N__10668\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5C_net\,
            ce => \N__10455\,
            sr => \N__10387\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10669\,
            in1 => \N__10544\,
            in2 => \_gnd_net_\,
            in3 => \N__10504\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10473\,
            ce => \N__10456\,
            sr => \N__10393\
        );

    \U712_BUFFERS.DRDDIR_i_m2_i_m2_LC_24_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001111111"
        )
    port map (
            in0 => \N__10270\,
            in1 => \N__10081\,
            in2 => \N__11103\,
            in3 => \N__10201\,
            lcout => \N_405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_DRDENn_0_a2_LC_24_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10082\,
            in1 => \N__11099\,
            in2 => \_gnd_net_\,
            in3 => \N__11074\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Sep 13 2025 21:18:14

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    ROM_DELAY : in std_logic_vector(1 downto 0);
    TM : in std_logic_vector(2 downto 0);
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : inout std_logic_vector(7 downto 4);
    RESETn : in std_logic;
    OVL : in std_logic;
    CONFIGENn : out std_logic;
    PPIO : out std_logic;
    PORTSIZE : out std_logic;
    TICK60 : out std_logic;
    PCS1 : out std_logic;
    CIACS0n : out std_logic;
    SCS0 : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    AGNUS_CLK : out std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    XCLK : in std_logic;
    CIACS1n : out std_logic;
    PPIO_J : in std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    PCS0 : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    XCLK_ENn : in std_logic;
    SCS1 : out std_logic;
    REGSPACEn : out std_logic;
    F_ENn : out std_logic;
    TSn : in std_logic;
    SPIO_J : in std_logic;
    SPIO : out std_logic;
    RTC_ENn : out std_logic;
    ATA_ENn : out std_logic;
    TACKn : inout std_logic;
    ROMENn : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__11620\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10825\ : std_logic;
signal \N__10822\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10762\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10753\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10738\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10688\ : std_logic;
signal \N__10685\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10663\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10652\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10592\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10577\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10571\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10544\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10538\ : std_logic;
signal \N__10535\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10434\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10390\ : std_logic;
signal \N__10387\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10363\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10122\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9958\ : std_logic;
signal \N__9953\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9947\ : std_logic;
signal \N__9946\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9794\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9791\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9788\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9753\ : std_logic;
signal \N__9750\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9585\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9518\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9405\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9282\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9273\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9213\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9056\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8987\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8921\ : std_logic;
signal \N__8918\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8912\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8906\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8637\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8446\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8387\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8330\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8312\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8267\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8227\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__8001\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7901\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7845\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7661\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7611\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7575\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7569\ : std_logic;
signal \N__7566\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7539\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7508\ : std_logic;
signal \N__7505\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7433\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7382\ : std_logic;
signal \N__7379\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7373\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7353\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7245\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7184\ : std_logic;
signal \N__7181\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7146\ : std_logic;
signal \N__7143\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7125\ : std_logic;
signal \N__7124\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7065\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7062\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7038\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6989\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6972\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6918\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6867\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6840\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6810\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6804\ : std_logic;
signal \N__6801\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6750\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6585\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6546\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6488\ : std_logic;
signal \N__6485\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6470\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6462\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6434\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5847\ : std_logic;
signal \N__5844\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5805\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5795\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5772\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5678\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5660\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5588\ : std_logic;
signal \N__5585\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5556\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5487\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5319\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5220\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5136\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5132\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5115\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5106\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4967\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4852\ : std_logic;
signal \N__4849\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4749\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4695\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4665\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4242\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4211\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \PPIO_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \SPIO_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_26\ : std_logic;
signal \A_c_25\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_29\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10\ : std_logic;
signal \N_61_i\ : std_logic;
signal \N_89_cascade_\ : std_logic;
signal \N_94_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \N_89\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8\ : std_logic;
signal \A_c_15\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_\ : std_logic;
signal \A_c_16\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \A_c_18\ : std_logic;
signal \A_c_17\ : std_logic;
signal \LIDE_BASE_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\ : std_logic;
signal \LIDE_BASE_4\ : std_logic;
signal \LIDE_BASE_3\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\ : std_logic;
signal \ATA_SPACE_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\ : std_logic;
signal \OVL_c\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE\ : std_logic;
signal \U409_ADDRESS_DECODE.N_34\ : std_logic;
signal \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4\ : std_logic;
signal \U409_AUTOCONFIG.N_227_3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.N_34_1\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0\ : std_logic;
signal \N_100\ : std_logic;
signal \N_94\ : std_logic;
signal \U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6_0_0\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_\ : std_logic;
signal \A_c_23\ : std_logic;
signal \U409_ADDRESS_DECODE.N_92\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_4\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_5\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \D_1_i\ : std_logic;
signal \D_in_4\ : std_logic;
signal \U409_AUTOCONFIG.N_76\ : std_logic;
signal \D_in_6\ : std_logic;
signal \D_in_5\ : std_logic;
signal \U409_AUTOCONFIG.N_82\ : std_logic;
signal \D_OUT_3\ : std_logic;
signal \U409_AUTOCONFIG.N_80\ : std_logic;
signal \LIDE_BASE_2\ : std_logic;
signal \LIDE_BASE_7\ : std_logic;
signal \U409_AUTOCONFIG.N_74\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\ : std_logic;
signal \A_c_22\ : std_logic;
signal \A_c_21\ : std_logic;
signal \LIDE_BASE_5\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.N_72\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6Z0Z_0\ : std_logic;
signal \LIDE_BASE_6\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_6C_net\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_0_2\ : std_logic;
signal \INVU409_AUTOCONFIG.PR_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_225\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_13Z0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_70\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\ : std_logic;
signal \D_OUT_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_BASE_10\ : std_logic;
signal \D_in_7\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_BASE_10_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_78\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_BASE_10_2\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_\ : std_logic;
signal \D_OUT_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_\ : std_logic;
signal \D_OUT_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1\ : std_logic;
signal \AUTOBOOT_c\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.N_214_0\ : std_logic;
signal \U409_AUTOCONFIG.N_193_1\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.N_159\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_192\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\ : std_logic;
signal \U409_AUTOCONFIG.N_184_0\ : std_logic;
signal \U409_AUTOCONFIG.N_167\ : std_logic;
signal \U409_AUTOCONFIG.N_213_i\ : std_logic;
signal \U409_AUTOCONFIG.N_182_0\ : std_logic;
signal \U409_AUTOCONFIG.N_223\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0\ : std_logic;
signal \A_c_3\ : std_logic;
signal \U409_AUTOCONFIG.N_190\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_1\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U409_AUTOCONFIG.N_198\ : std_logic;
signal \U409_AUTOCONFIG.N_222\ : std_logic;
signal \ATA_SPACE\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_AUTOCONFIG.D_OUT_sm0_0\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONFZ0\ : std_logic;
signal \INVU409_AUTOCONFIG.CONFIGENnC_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2\ : std_logic;
signal \U409_AUTOCONFIG.un1_AZ0Z_13\ : std_logic;
signal \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_0C_net\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \CONFIGURED\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_AUTOCONFIG.STATE4\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_1\ : std_logic;
signal \INVU409_AUTOCONFIG.AC_TACKC_net\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_TRANSFER_ACK.N_53\ : std_logic;
signal \U409_TRANSFER_ACK.N_53_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \TACK_OUT\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.N_62\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_CIA.CLK_CIA6_3_cascade_\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_2_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3\ : std_logic;
signal \U409_CIA.CLK_CIA6_0_cascade_\ : std_logic;
signal \U409_CIA.CLK_CIA6_3\ : std_logic;
signal \U409_CIA.CLK_CIA6_cascade_\ : std_logic;
signal \U409_CIA.CLK_CIA_RNOZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \TSn_c\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CLK_CIA6_0\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_19_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_23\ : std_logic;
signal \U409_TRANSFER_ACK.N_22\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENnC_net\ : std_logic;
signal \bfn_15_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_TRANSFER_ACK.N_101\ : std_logic;
signal \U409_TRANSFER_ACK.N_19\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\ : std_logic;
signal \ROMEN\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_11\ : std_logic;
signal \U409_TICK.TICK503_8_cascade_\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_8_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.TICK603_11\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.N_6_0\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_17_7_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \PCS1_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z0\ : std_logic;
signal \PCS0_c\ : std_logic;
signal \SCS0_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \SCS1_c\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \XCLK_c\ : std_logic;
signal \XCLK_ENn_c\ : std_logic;
signal \AGNUS_CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK6_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \CLK28_IN_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \SPIO_J_wire\ : std_logic;
signal \PPIO_wire\ : std_logic;
signal \PPIO_J_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AUTOBOOT_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \F_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \SCS1_wire\ : std_logic;
signal \AGNUS_CLK_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \XCLK_ENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \SPIO_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \PCS0_wire\ : std_logic;
signal \CLK_CIA_wire\ : std_logic;
signal \PCS1_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \SCS0_wire\ : std_logic;
signal \XCLK_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK6_wire\ <= CLK6;
    \CLK40_IN_wire\ <= CLK40_IN;
    \CLK28_IN_wire\ <= CLK28_IN;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \SPIO_J_wire\ <= SPIO_J;
    PPIO <= \PPIO_wire\;
    \PPIO_J_wire\ <= PPIO_J;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \AUTOBOOT_wire\ <= AUTOBOOT;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    F_ENn <= \F_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    SCS1 <= \SCS1_wire\;
    AGNUS_CLK <= \AGNUS_CLK_wire\;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \XCLK_ENn_wire\ <= XCLK_ENn;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    SPIO <= \SPIO_wire\;
    TICK60 <= \TICK60_wire\;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    PCS0 <= \PCS0_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    PCS1 <= \PCS1_wire\;
    BUFENn <= \BUFENn_wire\;
    SCS0 <= \SCS0_wire\;
    \XCLK_wire\ <= XCLK;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__7754\,
            RESETB => \N__10763\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11618\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11620\,
            DIN => \N__11619\,
            DOUT => \N__11618\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11620\,
            PADOUT => \N__11619\,
            PADIN => \N__11618\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11608\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11610\,
            DIN => \N__11609\,
            DOUT => \N__11608\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11610\,
            PADOUT => \N__11609\,
            PADIN => \N__11608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__11598\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11600\,
            DIN => \N__11599\,
            DOUT => \N__11598\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11600\,
            PADOUT => \N__11599\,
            PADIN => \N__11598\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11589\,
            DIN => \N__11588\,
            DOUT => \N__11587\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11589\,
            PADOUT => \N__11588\,
            PADIN => \N__11587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11580\,
            DIN => \N__11579\,
            DOUT => \N__11578\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11580\,
            PADOUT => \N__11579\,
            PADIN => \N__11578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11571\,
            DIN => \N__11570\,
            DOUT => \N__11569\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11571\,
            PADOUT => \N__11570\,
            PADIN => \N__11569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5510\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__5411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11562\,
            DIN => \N__11561\,
            DOUT => \N__11560\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11562\,
            PADOUT => \N__11561\,
            PADIN => \N__11560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11553\,
            DIN => \N__11552\,
            DOUT => \N__11551\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11553\,
            PADOUT => \N__11552\,
            PADIN => \N__11551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11544\,
            DIN => \N__11543\,
            DOUT => \N__11542\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11544\,
            PADOUT => \N__11543\,
            PADIN => \N__11542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4322\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11535\,
            DIN => \N__11534\,
            DOUT => \N__11533\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11535\,
            PADOUT => \N__11534\,
            PADIN => \N__11533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11526\,
            DIN => \N__11525\,
            DOUT => \N__11524\,
            PACKAGEPIN => \SPIO_J_wire\
        );

    \SPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11526\,
            PADOUT => \N__11525\,
            PADIN => \N__11524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11517\,
            DIN => \N__11516\,
            DOUT => \N__11515\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11517\,
            PADOUT => \N__11516\,
            PADIN => \N__11515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5487\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__6410\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11508\,
            DIN => \N__11507\,
            DOUT => \N__11506\,
            PACKAGEPIN => \PPIO_wire\
        );

    \PPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11508\,
            PADOUT => \N__11507\,
            PADIN => \N__11506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4271\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11499\,
            DIN => \N__11498\,
            DOUT => \N__11497\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11499\,
            PADOUT => \N__11498\,
            PADIN => \N__11497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11490\,
            DIN => \N__11489\,
            DOUT => \N__11488\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11490\,
            PADOUT => \N__11489\,
            PADIN => \N__11488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11481\,
            DIN => \N__11480\,
            DOUT => \N__11479\,
            PACKAGEPIN => \PPIO_J_wire\
        );

    \PPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11481\,
            PADOUT => \N__11480\,
            PADIN => \N__11479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11472\,
            DIN => \N__11471\,
            DOUT => \N__11470\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11472\,
            PADOUT => \N__11471\,
            PADIN => \N__11470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4772\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11463\,
            DIN => \N__11462\,
            DOUT => \N__11461\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11463\,
            PADOUT => \N__11462\,
            PADIN => \N__11461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11454\,
            DIN => \N__11453\,
            DOUT => \N__11452\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11454\,
            PADOUT => \N__11453\,
            PADIN => \N__11452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11445\,
            DIN => \N__11444\,
            DOUT => \N__11443\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11445\,
            PADOUT => \N__11444\,
            PADIN => \N__11443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9137\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AUTOBOOT_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__11436\,
            DIN => \N__11435\,
            DOUT => \N__11434\,
            PACKAGEPIN => \AUTOBOOT_wire\
        );

    \AUTOBOOT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11436\,
            PADOUT => \N__11435\,
            PADIN => \N__11434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AUTOBOOT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11427\,
            DIN => \N__11426\,
            DOUT => \N__11425\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11427\,
            PADOUT => \N__11426\,
            PADIN => \N__11425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11418\,
            DIN => \N__11417\,
            DOUT => \N__11416\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11418\,
            PADOUT => \N__11417\,
            PADIN => \N__11416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5303\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11409\,
            DIN => \N__11408\,
            DOUT => \N__11407\,
            PACKAGEPIN => \F_ENn_wire\
        );

    \F_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11409\,
            PADOUT => \N__11408\,
            PADIN => \N__11407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10762\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11400\,
            DIN => \N__11399\,
            DOUT => \N__11398\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11400\,
            PADOUT => \N__11399\,
            PADIN => \N__11398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11391\,
            DIN => \N__11390\,
            DOUT => \N__11389\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11391\,
            PADOUT => \N__11390\,
            PADIN => \N__11389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11382\,
            DIN => \N__11381\,
            DOUT => \N__11380\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11382\,
            PADOUT => \N__11381\,
            PADIN => \N__11380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11373\,
            DIN => \N__11372\,
            DOUT => \N__11371\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11373\,
            PADOUT => \N__11372\,
            PADIN => \N__11371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11364\,
            DIN => \N__11363\,
            DOUT => \N__11362\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11364\,
            PADOUT => \N__11363\,
            PADIN => \N__11362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11355\,
            DIN => \N__11354\,
            DOUT => \N__11353\,
            PACKAGEPIN => \SCS1_wire\
        );

    \SCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11355\,
            PADOUT => \N__11354\,
            PADIN => \N__11353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10928\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11346\,
            DIN => \N__11345\,
            DOUT => \N__11344\,
            PACKAGEPIN => \AGNUS_CLK_wire\
        );

    \AGNUS_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11346\,
            PADOUT => \N__11345\,
            PADIN => \N__11344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10865\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11337\,
            DIN => \N__11336\,
            DOUT => \N__11335\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11337\,
            PADOUT => \N__11336\,
            PADIN => \N__11335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11328\,
            DIN => \N__11327\,
            DOUT => \N__11326\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11328\,
            PADOUT => \N__11327\,
            PADIN => \N__11326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11319\,
            DIN => \N__11318\,
            DOUT => \N__11317\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11319\,
            PADOUT => \N__11318\,
            PADIN => \N__11317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9062\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11310\,
            DIN => \N__11309\,
            DOUT => \N__11308\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11310\,
            PADOUT => \N__11309\,
            PADIN => \N__11308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11301\,
            DIN => \N__11300\,
            DOUT => \N__11299\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11301\,
            PADOUT => \N__11300\,
            PADIN => \N__11299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11292\,
            DIN => \N__11291\,
            DOUT => \N__11290\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11292\,
            PADOUT => \N__11291\,
            PADIN => \N__11290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11283\,
            DIN => \N__11282\,
            DOUT => \N__11281\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11283\,
            PADOUT => \N__11282\,
            PADIN => \N__11281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11274\,
            DIN => \N__11273\,
            DOUT => \N__11272\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11274\,
            PADOUT => \N__11273\,
            PADIN => \N__11272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9083\,
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11265\,
            DIN => \N__11264\,
            DOUT => \N__11263\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11265\,
            PADOUT => \N__11264\,
            PADIN => \N__11263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5505\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__6056\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11256\,
            DIN => \N__11255\,
            DOUT => \N__11254\,
            PACKAGEPIN => \XCLK_ENn_wire\
        );

    \XCLK_ENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11256\,
            PADOUT => \N__11255\,
            PADIN => \N__11254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_ENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11247\,
            DIN => \N__11246\,
            DOUT => \N__11245\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11247\,
            PADOUT => \N__11246\,
            PADIN => \N__11245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11238\,
            DIN => \N__11237\,
            DOUT => \N__11236\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11238\,
            PADOUT => \N__11237\,
            PADIN => \N__11236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11229\,
            DIN => \N__11228\,
            DOUT => \N__11227\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11229\,
            PADOUT => \N__11228\,
            PADIN => \N__11227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11220\,
            DIN => \N__11219\,
            DOUT => \N__11218\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11220\,
            PADOUT => \N__11219\,
            PADIN => \N__11218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7328\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11211\,
            DIN => \N__11210\,
            DOUT => \N__11209\,
            PACKAGEPIN => \SPIO_wire\
        );

    \SPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11211\,
            PADOUT => \N__11210\,
            PADIN => \N__11209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4307\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11202\,
            DIN => \N__11201\,
            DOUT => \N__11200\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11202\,
            PADOUT => \N__11201\,
            PADIN => \N__11200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9557\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11193\,
            DIN => \N__11192\,
            DOUT => \N__11191\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11193\,
            PADOUT => \N__11192\,
            PADIN => \N__11191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11184\,
            DIN => \N__11183\,
            DOUT => \N__11182\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11184\,
            PADOUT => \N__11183\,
            PADIN => \N__11182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11175\,
            DIN => \N__11174\,
            DOUT => \N__11173\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11175\,
            PADOUT => \N__11174\,
            PADIN => \N__11173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11166\,
            DIN => \N__11165\,
            DOUT => \N__11164\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11166\,
            PADOUT => \N__11165\,
            PADIN => \N__11164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10700\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11157\,
            DIN => \N__11156\,
            DOUT => \N__11155\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11157\,
            PADOUT => \N__11156\,
            PADIN => \N__11155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11148\,
            DIN => \N__11147\,
            DOUT => \N__11146\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11148\,
            PADOUT => \N__11147\,
            PADIN => \N__11146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8435\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11139\,
            DIN => \N__11138\,
            DOUT => \N__11137\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11139\,
            PADOUT => \N__11138\,
            PADIN => \N__11137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5534\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11130\,
            DIN => \N__11129\,
            DOUT => \N__11128\,
            PACKAGEPIN => \PCS0_wire\
        );

    \PCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11130\,
            PADOUT => \N__11129\,
            PADIN => \N__11128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10649\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11121\,
            DIN => \N__11120\,
            DOUT => \N__11119\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11121\,
            PADOUT => \N__11120\,
            PADIN => \N__11119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11112\,
            DIN => \N__11111\,
            DOUT => \N__11110\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11112\,
            PADOUT => \N__11111\,
            PADIN => \N__11110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8918\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11103\,
            DIN => \N__11102\,
            DOUT => \N__11101\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11103\,
            PADOUT => \N__11102\,
            PADIN => \N__11101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11094\,
            DIN => \N__11093\,
            DOUT => \N__11092\,
            PACKAGEPIN => \PCS1_wire\
        );

    \PCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11094\,
            PADOUT => \N__11093\,
            PADIN => \N__11092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10691\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11085\,
            DIN => \N__11084\,
            DOUT => \N__11083\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11085\,
            PADOUT => \N__11084\,
            PADIN => \N__11083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9133\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__8159\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11076\,
            DIN => \N__11075\,
            DOUT => \N__11074\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11076\,
            PADOUT => \N__11075\,
            PADIN => \N__11074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11067\,
            DIN => \N__11066\,
            DOUT => \N__11065\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11067\,
            PADOUT => \N__11066\,
            PADIN => \N__11065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7382\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11058\,
            DIN => \N__11057\,
            DOUT => \N__11056\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11058\,
            PADOUT => \N__11057\,
            PADIN => \N__11056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11049\,
            DIN => \N__11048\,
            DOUT => \N__11047\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11049\,
            PADOUT => \N__11048\,
            PADIN => \N__11047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5506\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__6194\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11040\,
            DIN => \N__11039\,
            DOUT => \N__11038\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11040\,
            PADOUT => \N__11039\,
            PADIN => \N__11038\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11031\,
            DIN => \N__11030\,
            DOUT => \N__11029\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11031\,
            PADOUT => \N__11030\,
            PADIN => \N__11029\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11022\,
            DIN => \N__11021\,
            DOUT => \N__11020\,
            PACKAGEPIN => \SCS0_wire\
        );

    \SCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11022\,
            PADOUT => \N__11021\,
            PADIN => \N__11020\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10634\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11013\,
            DIN => \N__11012\,
            DOUT => \N__11011\,
            PACKAGEPIN => \XCLK_wire\
        );

    \XCLK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11013\,
            PADOUT => \N__11012\,
            PADIN => \N__11011\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11004\,
            DIN => \N__11003\,
            DOUT => \N__11002\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11004\,
            PADOUT => \N__11003\,
            PADIN => \N__11002\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__10995\,
            DIN => \N__10994\,
            DOUT => \N__10993\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__10995\,
            PADOUT => \N__10994\,
            PADIN => \N__10993\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2625\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10970\
        );

    \I__2624\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10970\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10967\
        );

    \I__2622\ : Sp12to4
    port map (
            O => \N__10967\,
            I => \N__10964\
        );

    \I__2621\ : Span12Mux_h
    port map (
            O => \N__10964\,
            I => \N__10961\
        );

    \I__2620\ : Odrv12
    port map (
            O => \N__10961\,
            I => \U409_ADDRESS_DECODE.CSZ0Z1\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10948\
        );

    \I__2618\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10948\
        );

    \I__2617\ : InMux
    port map (
            O => \N__10956\,
            I => \N__10948\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10955\,
            I => \N__10945\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10940\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__10945\,
            I => \N__10940\
        );

    \I__2613\ : Span12Mux_v
    port map (
            O => \N__10940\,
            I => \N__10937\
        );

    \I__2612\ : Span12Mux_h
    port map (
            O => \N__10937\,
            I => \N__10934\
        );

    \I__2611\ : Span12Mux_h
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__2610\ : Odrv12
    port map (
            O => \N__10931\,
            I => \A_c_14\
        );

    \I__2609\ : IoInMux
    port map (
            O => \N__10928\,
            I => \N__10925\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__2607\ : Span12Mux_s4_h
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__2606\ : Odrv12
    port map (
            O => \N__10919\,
            I => \SCS1_c\
        );

    \I__2605\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__10913\,
            I => \N__10906\
        );

    \I__2603\ : ClkMux
    port map (
            O => \N__10912\,
            I => \N__10895\
        );

    \I__2602\ : ClkMux
    port map (
            O => \N__10911\,
            I => \N__10895\
        );

    \I__2601\ : ClkMux
    port map (
            O => \N__10910\,
            I => \N__10895\
        );

    \I__2600\ : ClkMux
    port map (
            O => \N__10909\,
            I => \N__10895\
        );

    \I__2599\ : Glb2LocalMux
    port map (
            O => \N__10906\,
            I => \N__10895\
        );

    \I__2598\ : GlobalMux
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__2597\ : gio2CtrlBuf
    port map (
            O => \N__10892\,
            I => \CLK28_IN_c_g\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__2593\ : Odrv4
    port map (
            O => \N__10880\,
            I => \XCLK_c\
        );

    \I__2592\ : InMux
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__10874\,
            I => \N__10871\
        );

    \I__2590\ : Span12Mux_v
    port map (
            O => \N__10871\,
            I => \N__10868\
        );

    \I__2589\ : Odrv12
    port map (
            O => \N__10868\,
            I => \XCLK_ENn_c\
        );

    \I__2588\ : IoInMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10859\
        );

    \I__2586\ : Span4Mux_s3_h
    port map (
            O => \N__10859\,
            I => \N__10856\
        );

    \I__2585\ : Odrv4
    port map (
            O => \N__10856\,
            I => \AGNUS_CLK_c\
        );

    \I__2584\ : InMux
    port map (
            O => \N__10853\,
            I => \N__10849\
        );

    \I__2583\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10846\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__10849\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__10846\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__2579\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10835\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__2577\ : InMux
    port map (
            O => \N__10832\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__2576\ : InMux
    port map (
            O => \N__10829\,
            I => \N__10825\
        );

    \I__2575\ : InMux
    port map (
            O => \N__10828\,
            I => \N__10822\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__10825\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2573\ : LocalMux
    port map (
            O => \N__10822\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10817\,
            I => \N__10814\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__10814\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__2570\ : InMux
    port map (
            O => \N__10811\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__2569\ : InMux
    port map (
            O => \N__10808\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10801\
        );

    \I__2567\ : InMux
    port map (
            O => \N__10804\,
            I => \N__10798\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__10801\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__10798\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__2564\ : ClkMux
    port map (
            O => \N__10793\,
            I => \N__10769\
        );

    \I__2563\ : ClkMux
    port map (
            O => \N__10792\,
            I => \N__10769\
        );

    \I__2562\ : ClkMux
    port map (
            O => \N__10791\,
            I => \N__10769\
        );

    \I__2561\ : ClkMux
    port map (
            O => \N__10790\,
            I => \N__10769\
        );

    \I__2560\ : ClkMux
    port map (
            O => \N__10789\,
            I => \N__10769\
        );

    \I__2559\ : ClkMux
    port map (
            O => \N__10788\,
            I => \N__10769\
        );

    \I__2558\ : ClkMux
    port map (
            O => \N__10787\,
            I => \N__10769\
        );

    \I__2557\ : ClkMux
    port map (
            O => \N__10786\,
            I => \N__10769\
        );

    \I__2556\ : GlobalMux
    port map (
            O => \N__10769\,
            I => \N__10766\
        );

    \I__2555\ : gio2CtrlBuf
    port map (
            O => \N__10766\,
            I => \CLK6_c_g\
        );

    \I__2554\ : IoInMux
    port map (
            O => \N__10763\,
            I => \N__10759\
        );

    \I__2553\ : IoInMux
    port map (
            O => \N__10762\,
            I => \N__10756\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10759\,
            I => \N__10753\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__10756\,
            I => \N__10750\
        );

    \I__2550\ : IoSpan4Mux
    port map (
            O => \N__10753\,
            I => \N__10747\
        );

    \I__2549\ : IoSpan4Mux
    port map (
            O => \N__10750\,
            I => \N__10744\
        );

    \I__2548\ : Sp12to4
    port map (
            O => \N__10747\,
            I => \N__10741\
        );

    \I__2547\ : Span4Mux_s2_h
    port map (
            O => \N__10744\,
            I => \N__10738\
        );

    \I__2546\ : Span12Mux_s9_v
    port map (
            O => \N__10741\,
            I => \N__10735\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__10738\,
            I => \N__10732\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__10735\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2543\ : Odrv4
    port map (
            O => \N__10732\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10727\,
            I => \N__10724\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__10724\,
            I => \N__10721\
        );

    \I__2540\ : Span4Mux_v
    port map (
            O => \N__10721\,
            I => \N__10718\
        );

    \I__2539\ : Span4Mux_h
    port map (
            O => \N__10718\,
            I => \N__10714\
        );

    \I__2538\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10711\
        );

    \I__2537\ : Sp12to4
    port map (
            O => \N__10714\,
            I => \N__10708\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10705\
        );

    \I__2535\ : Odrv12
    port map (
            O => \N__10708\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__10705\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn\
        );

    \I__2533\ : IoInMux
    port map (
            O => \N__10700\,
            I => \N__10697\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2531\ : Odrv12
    port map (
            O => \N__10694\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__2530\ : IoInMux
    port map (
            O => \N__10691\,
            I => \N__10688\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10688\,
            I => \N__10685\
        );

    \I__2528\ : IoSpan4Mux
    port map (
            O => \N__10685\,
            I => \N__10682\
        );

    \I__2527\ : Span4Mux_s3_h
    port map (
            O => \N__10682\,
            I => \N__10679\
        );

    \I__2526\ : Odrv4
    port map (
            O => \N__10679\,
            I => \PCS1_c\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10676\,
            I => \N__10673\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__10673\,
            I => \N__10669\
        );

    \I__2523\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10666\
        );

    \I__2522\ : Sp12to4
    port map (
            O => \N__10669\,
            I => \N__10663\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10666\,
            I => \N__10660\
        );

    \I__2520\ : Span12Mux_v
    port map (
            O => \N__10663\,
            I => \N__10655\
        );

    \I__2519\ : Sp12to4
    port map (
            O => \N__10660\,
            I => \N__10655\
        );

    \I__2518\ : Span12Mux_h
    port map (
            O => \N__10655\,
            I => \N__10652\
        );

    \I__2517\ : Odrv12
    port map (
            O => \N__10652\,
            I => \U409_ADDRESS_DECODE.CSZ0Z0\
        );

    \I__2516\ : IoInMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__2514\ : Span4Mux_s3_h
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__2513\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__2512\ : Odrv4
    port map (
            O => \N__10637\,
            I => \PCS0_c\
        );

    \I__2511\ : IoInMux
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10631\,
            I => \N__10628\
        );

    \I__2509\ : Span4Mux_s3_h
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__10622\,
            I => \SCS0_c\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__10619\,
            I => \N__10616\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10612\
        );

    \I__2504\ : InMux
    port map (
            O => \N__10615\,
            I => \N__10609\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10612\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2502\ : LocalMux
    port map (
            O => \N__10609\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__10604\,
            I => \N__10601\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10598\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10598\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2498\ : InMux
    port map (
            O => \N__10595\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__10592\,
            I => \N__10589\
        );

    \I__2496\ : InMux
    port map (
            O => \N__10589\,
            I => \N__10585\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10582\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__10585\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__10582\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10577\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2491\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10571\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10571\,
            I => \N__10567\
        );

    \I__2489\ : InMux
    port map (
            O => \N__10570\,
            I => \N__10564\
        );

    \I__2488\ : Odrv4
    port map (
            O => \N__10567\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__10564\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2486\ : InMux
    port map (
            O => \N__10559\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2485\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10552\
        );

    \I__2484\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10549\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10552\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10549\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2481\ : InMux
    port map (
            O => \N__10544\,
            I => \N__10541\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10541\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10538\,
            I => \bfn_17_7_0_\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10535\,
            I => \N__10531\
        );

    \I__2477\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10528\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10531\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__10528\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10523\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10516\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10519\,
            I => \N__10513\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__10516\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10513\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__2469\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10505\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10505\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__2467\ : InMux
    port map (
            O => \N__10502\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2466\ : InMux
    port map (
            O => \N__10499\,
            I => \N__10495\
        );

    \I__2465\ : InMux
    port map (
            O => \N__10498\,
            I => \N__10492\
        );

    \I__2464\ : LocalMux
    port map (
            O => \N__10495\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10492\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10487\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2461\ : InMux
    port map (
            O => \N__10484\,
            I => \N__10480\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10477\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10480\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10477\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10472\,
            I => \N__10469\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10469\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10466\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10463\,
            I => \N__10458\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10462\,
            I => \N__10453\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10453\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10458\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10453\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10442\
        );

    \I__2448\ : InMux
    port map (
            O => \N__10447\,
            I => \N__10442\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10442\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10436\,
            I => \N__10427\
        );

    \I__2444\ : InMux
    port map (
            O => \N__10435\,
            I => \N__10427\
        );

    \I__2443\ : InMux
    port map (
            O => \N__10434\,
            I => \N__10427\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10427\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10421\,
            I => \N__10414\
        );

    \I__2439\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10414\
        );

    \I__2438\ : CascadeMux
    port map (
            O => \N__10419\,
            I => \N__10409\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__10414\,
            I => \N__10399\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10413\,
            I => \N__10395\
        );

    \I__2435\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10390\
        );

    \I__2434\ : InMux
    port map (
            O => \N__10409\,
            I => \N__10387\
        );

    \I__2433\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10384\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__10407\,
            I => \N__10381\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__10406\,
            I => \N__10378\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__10405\,
            I => \N__10371\
        );

    \I__2429\ : CascadeMux
    port map (
            O => \N__10404\,
            I => \N__10368\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__10403\,
            I => \N__10365\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__10402\,
            I => \N__10358\
        );

    \I__2426\ : Span4Mux_h
    port map (
            O => \N__10399\,
            I => \N__10355\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10352\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10395\,
            I => \N__10349\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10346\
        );

    \I__2422\ : InMux
    port map (
            O => \N__10393\,
            I => \N__10343\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10390\,
            I => \N__10340\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10387\,
            I => \N__10337\
        );

    \I__2419\ : InMux
    port map (
            O => \N__10384\,
            I => \N__10334\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10381\,
            I => \N__10329\
        );

    \I__2417\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10329\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10326\
        );

    \I__2415\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10323\
        );

    \I__2414\ : InMux
    port map (
            O => \N__10375\,
            I => \N__10318\
        );

    \I__2413\ : InMux
    port map (
            O => \N__10374\,
            I => \N__10318\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10315\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10306\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10365\,
            I => \N__10306\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10364\,
            I => \N__10306\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10363\,
            I => \N__10306\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__10362\,
            I => \N__10302\
        );

    \I__2406\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10297\
        );

    \I__2405\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10297\
        );

    \I__2404\ : Span4Mux_h
    port map (
            O => \N__10355\,
            I => \N__10294\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10352\,
            I => \N__10291\
        );

    \I__2402\ : Span4Mux_v
    port map (
            O => \N__10349\,
            I => \N__10287\
        );

    \I__2401\ : LocalMux
    port map (
            O => \N__10346\,
            I => \N__10284\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__10343\,
            I => \N__10281\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__10340\,
            I => \N__10272\
        );

    \I__2398\ : Span4Mux_v
    port map (
            O => \N__10337\,
            I => \N__10272\
        );

    \I__2397\ : LocalMux
    port map (
            O => \N__10334\,
            I => \N__10272\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10329\,
            I => \N__10272\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10326\,
            I => \N__10260\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__10323\,
            I => \N__10260\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10260\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__10315\,
            I => \N__10260\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10306\,
            I => \N__10260\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10305\,
            I => \N__10255\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10255\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10297\,
            I => \N__10252\
        );

    \I__2387\ : Span4Mux_h
    port map (
            O => \N__10294\,
            I => \N__10247\
        );

    \I__2386\ : Span4Mux_v
    port map (
            O => \N__10291\,
            I => \N__10247\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10244\
        );

    \I__2384\ : Span4Mux_v
    port map (
            O => \N__10287\,
            I => \N__10239\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__10284\,
            I => \N__10239\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10281\,
            I => \N__10234\
        );

    \I__2381\ : Span4Mux_v
    port map (
            O => \N__10272\,
            I => \N__10234\
        );

    \I__2380\ : InMux
    port map (
            O => \N__10271\,
            I => \N__10231\
        );

    \I__2379\ : Span4Mux_v
    port map (
            O => \N__10260\,
            I => \N__10228\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10255\,
            I => \N__10225\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10252\,
            I => \N__10218\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__10247\,
            I => \N__10218\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10244\,
            I => \N__10218\
        );

    \I__2374\ : Span4Mux_h
    port map (
            O => \N__10239\,
            I => \N__10215\
        );

    \I__2373\ : Span4Mux_h
    port map (
            O => \N__10234\,
            I => \N__10212\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10209\
        );

    \I__2371\ : Span4Mux_h
    port map (
            O => \N__10228\,
            I => \N__10204\
        );

    \I__2370\ : Span4Mux_v
    port map (
            O => \N__10225\,
            I => \N__10204\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__10218\,
            I => \N__10201\
        );

    \I__2368\ : Sp12to4
    port map (
            O => \N__10215\,
            I => \N__10196\
        );

    \I__2367\ : Sp12to4
    port map (
            O => \N__10212\,
            I => \N__10196\
        );

    \I__2366\ : Span12Mux_v
    port map (
            O => \N__10209\,
            I => \N__10189\
        );

    \I__2365\ : Sp12to4
    port map (
            O => \N__10204\,
            I => \N__10189\
        );

    \I__2364\ : Sp12to4
    port map (
            O => \N__10201\,
            I => \N__10189\
        );

    \I__2363\ : Span12Mux_h
    port map (
            O => \N__10196\,
            I => \N__10186\
        );

    \I__2362\ : Span12Mux_v
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__2361\ : Span12Mux_v
    port map (
            O => \N__10186\,
            I => \N__10178\
        );

    \I__2360\ : Span12Mux_h
    port map (
            O => \N__10183\,
            I => \N__10178\
        );

    \I__2359\ : Odrv12
    port map (
            O => \N__10178\,
            I => \RESETn_c\
        );

    \I__2358\ : InMux
    port map (
            O => \N__10175\,
            I => \N__10172\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10168\
        );

    \I__2356\ : InMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10168\,
            I => \N__10161\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10165\,
            I => \N__10158\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10155\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__10161\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__10158\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10155\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10148\,
            I => \N__10142\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10147\,
            I => \N__10135\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10135\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10145\,
            I => \N__10135\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10142\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10135\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2343\ : SRMux
    port map (
            O => \N__10130\,
            I => \N__10097\
        );

    \I__2342\ : SRMux
    port map (
            O => \N__10129\,
            I => \N__10097\
        );

    \I__2341\ : SRMux
    port map (
            O => \N__10128\,
            I => \N__10097\
        );

    \I__2340\ : SRMux
    port map (
            O => \N__10127\,
            I => \N__10097\
        );

    \I__2339\ : SRMux
    port map (
            O => \N__10126\,
            I => \N__10097\
        );

    \I__2338\ : SRMux
    port map (
            O => \N__10125\,
            I => \N__10097\
        );

    \I__2337\ : SRMux
    port map (
            O => \N__10124\,
            I => \N__10097\
        );

    \I__2336\ : SRMux
    port map (
            O => \N__10123\,
            I => \N__10097\
        );

    \I__2335\ : SRMux
    port map (
            O => \N__10122\,
            I => \N__10097\
        );

    \I__2334\ : SRMux
    port map (
            O => \N__10121\,
            I => \N__10097\
        );

    \I__2333\ : SRMux
    port map (
            O => \N__10120\,
            I => \N__10097\
        );

    \I__2332\ : GlobalMux
    port map (
            O => \N__10097\,
            I => \N__10094\
        );

    \I__2331\ : gio2CtrlBuf
    port map (
            O => \N__10094\,
            I => \RESETn_c_i_g\
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__10091\,
            I => \N__10087\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10084\
        );

    \I__2328\ : InMux
    port map (
            O => \N__10087\,
            I => \N__10078\
        );

    \I__2327\ : InMux
    port map (
            O => \N__10084\,
            I => \N__10078\
        );

    \I__2326\ : InMux
    port map (
            O => \N__10083\,
            I => \N__10075\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__10078\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__10075\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__10070\,
            I => \N__10066\
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__10069\,
            I => \N__10061\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10066\,
            I => \N__10058\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10065\,
            I => \N__10053\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10053\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10050\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__10058\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__10053\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10050\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2314\ : InMux
    port map (
            O => \N__10043\,
            I => \N__10039\
        );

    \I__2313\ : InMux
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__10039\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__10036\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2310\ : InMux
    port map (
            O => \N__10031\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10028\,
            I => \N__10024\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10024\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10021\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10016\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2304\ : InMux
    port map (
            O => \N__10013\,
            I => \N__10009\
        );

    \I__2303\ : InMux
    port map (
            O => \N__10012\,
            I => \N__10006\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10009\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10006\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2300\ : InMux
    port map (
            O => \N__10001\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9998\,
            I => \N__9994\
        );

    \I__2298\ : InMux
    port map (
            O => \N__9997\,
            I => \N__9991\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9994\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9991\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2295\ : CascadeMux
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__2294\ : InMux
    port map (
            O => \N__9983\,
            I => \N__9980\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9980\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9977\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__9974\,
            I => \N__9971\
        );

    \I__2290\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9968\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9968\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2288\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9961\
        );

    \I__2287\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9958\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__9961\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2285\ : LocalMux
    port map (
            O => \N__9958\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2284\ : InMux
    port map (
            O => \N__9953\,
            I => \N__9950\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9950\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9947\,
            I => \N__9943\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9946\,
            I => \N__9940\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__9943\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9940\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2278\ : CascadeMux
    port map (
            O => \N__9935\,
            I => \N__9928\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__9934\,
            I => \N__9924\
        );

    \I__2276\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9921\
        );

    \I__2275\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9918\
        );

    \I__2274\ : InMux
    port map (
            O => \N__9931\,
            I => \N__9915\
        );

    \I__2273\ : InMux
    port map (
            O => \N__9928\,
            I => \N__9912\
        );

    \I__2272\ : InMux
    port map (
            O => \N__9927\,
            I => \N__9909\
        );

    \I__2271\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9906\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__9921\,
            I => \N__9900\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__9918\,
            I => \N__9892\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__9915\,
            I => \N__9886\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__9912\,
            I => \N__9883\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__9909\,
            I => \N__9880\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__9906\,
            I => \N__9877\
        );

    \I__2264\ : ClkMux
    port map (
            O => \N__9905\,
            I => \N__9842\
        );

    \I__2263\ : ClkMux
    port map (
            O => \N__9904\,
            I => \N__9842\
        );

    \I__2262\ : ClkMux
    port map (
            O => \N__9903\,
            I => \N__9842\
        );

    \I__2261\ : Glb2LocalMux
    port map (
            O => \N__9900\,
            I => \N__9842\
        );

    \I__2260\ : ClkMux
    port map (
            O => \N__9899\,
            I => \N__9842\
        );

    \I__2259\ : ClkMux
    port map (
            O => \N__9898\,
            I => \N__9842\
        );

    \I__2258\ : ClkMux
    port map (
            O => \N__9897\,
            I => \N__9842\
        );

    \I__2257\ : ClkMux
    port map (
            O => \N__9896\,
            I => \N__9842\
        );

    \I__2256\ : ClkMux
    port map (
            O => \N__9895\,
            I => \N__9842\
        );

    \I__2255\ : Glb2LocalMux
    port map (
            O => \N__9892\,
            I => \N__9842\
        );

    \I__2254\ : ClkMux
    port map (
            O => \N__9891\,
            I => \N__9842\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9890\,
            I => \N__9842\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9889\,
            I => \N__9842\
        );

    \I__2251\ : Glb2LocalMux
    port map (
            O => \N__9886\,
            I => \N__9842\
        );

    \I__2250\ : Glb2LocalMux
    port map (
            O => \N__9883\,
            I => \N__9842\
        );

    \I__2249\ : Glb2LocalMux
    port map (
            O => \N__9880\,
            I => \N__9842\
        );

    \I__2248\ : Glb2LocalMux
    port map (
            O => \N__9877\,
            I => \N__9842\
        );

    \I__2247\ : GlobalMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__2246\ : gio2CtrlBuf
    port map (
            O => \N__9839\,
            I => \CLK40_IN_c_g\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9833\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__9833\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2243\ : CascadeMux
    port map (
            O => \N__9830\,
            I => \U409_TRANSFER_ACK.N_17_mux_cascade_\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__9824\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\
        );

    \I__2240\ : CascadeMux
    port map (
            O => \N__9821\,
            I => \U409_TRANSFER_ACK.N_3_0_cascade_\
        );

    \I__2239\ : InMux
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__9815\,
            I => \U409_TRANSFER_ACK.N_6_0\
        );

    \I__2237\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9809\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2235\ : InMux
    port map (
            O => \N__9806\,
            I => \N__9802\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9805\,
            I => \N__9799\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__9802\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9799\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2231\ : InMux
    port map (
            O => \N__9794\,
            I => \N__9781\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9793\,
            I => \N__9781\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9792\,
            I => \N__9781\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9791\,
            I => \N__9772\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9790\,
            I => \N__9772\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9772\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9788\,
            I => \N__9772\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__9781\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__9772\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2222\ : CascadeMux
    port map (
            O => \N__9767\,
            I => \N__9760\
        );

    \I__2221\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \N__9757\
        );

    \I__2220\ : CascadeMux
    port map (
            O => \N__9765\,
            I => \N__9754\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__9764\,
            I => \N__9750\
        );

    \I__2218\ : InMux
    port map (
            O => \N__9763\,
            I => \N__9737\
        );

    \I__2217\ : InMux
    port map (
            O => \N__9760\,
            I => \N__9737\
        );

    \I__2216\ : InMux
    port map (
            O => \N__9757\,
            I => \N__9737\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9737\
        );

    \I__2214\ : InMux
    port map (
            O => \N__9753\,
            I => \N__9737\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9750\,
            I => \N__9730\
        );

    \I__2212\ : InMux
    port map (
            O => \N__9749\,
            I => \N__9730\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9730\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9737\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__9730\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__9725\,
            I => \N__9721\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__9724\,
            I => \N__9717\
        );

    \I__2206\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9705\
        );

    \I__2205\ : InMux
    port map (
            O => \N__9720\,
            I => \N__9705\
        );

    \I__2204\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9705\
        );

    \I__2203\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9694\
        );

    \I__2202\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9694\
        );

    \I__2201\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9694\
        );

    \I__2200\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9694\
        );

    \I__2199\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9694\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__9705\,
            I => \N__9691\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9694\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2196\ : Odrv4
    port map (
            O => \N__9691\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2195\ : InMux
    port map (
            O => \N__9686\,
            I => \N__9683\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__9683\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2193\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9676\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__9676\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9673\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9662\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__9662\,
            I => \N__9655\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9652\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9645\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9659\,
            I => \N__9645\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9658\,
            I => \N__9645\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__9655\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9652\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__9645\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2179\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__9635\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__2177\ : InMux
    port map (
            O => \N__9632\,
            I => \N__9629\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__9629\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__9626\,
            I => \N__9620\
        );

    \I__2174\ : InMux
    port map (
            O => \N__9625\,
            I => \N__9607\
        );

    \I__2173\ : InMux
    port map (
            O => \N__9624\,
            I => \N__9607\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9607\
        );

    \I__2171\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9607\
        );

    \I__2170\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9598\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9618\,
            I => \N__9598\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9598\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9598\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9607\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__9598\,
            I => \U409_TICK.TICK503_10\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9574\
        );

    \I__2163\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9574\
        );

    \I__2162\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9574\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9574\
        );

    \I__2160\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9574\
        );

    \I__2159\ : InMux
    port map (
            O => \N__9588\,
            I => \N__9565\
        );

    \I__2158\ : InMux
    port map (
            O => \N__9587\,
            I => \N__9565\
        );

    \I__2157\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9565\
        );

    \I__2156\ : InMux
    port map (
            O => \N__9585\,
            I => \N__9565\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__9574\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9565\,
            I => \U409_TICK.TICK503_14\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__9560\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2152\ : IoInMux
    port map (
            O => \N__9557\,
            I => \N__9554\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__2150\ : Span4Mux_s1_v
    port map (
            O => \N__9551\,
            I => \N__9548\
        );

    \I__2149\ : Sp12to4
    port map (
            O => \N__9548\,
            I => \N__9545\
        );

    \I__2148\ : Span12Mux_h
    port map (
            O => \N__9545\,
            I => \N__9541\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9544\,
            I => \N__9538\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__9541\,
            I => \TICK60_c\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__9538\,
            I => \TICK60_c\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9533\,
            I => \N__9529\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9529\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9526\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2140\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9518\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9518\,
            I => \N__9514\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9517\,
            I => \N__9511\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__9514\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9511\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__9506\,
            I => \U409_TICK.TICK603_8_cascade_\
        );

    \I__2134\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9499\
        );

    \I__2133\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9496\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__9499\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9496\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__9491\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__2129\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9484\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__9487\,
            I => \N__9479\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__9484\,
            I => \N__9476\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9483\,
            I => \N__9473\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9470\
        );

    \I__2124\ : InMux
    port map (
            O => \N__9479\,
            I => \N__9467\
        );

    \I__2123\ : Odrv4
    port map (
            O => \N__9476\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9473\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__9470\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9467\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2119\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9455\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__9455\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__9452\,
            I => \N__9449\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9446\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__9446\,
            I => \N__9442\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__2113\ : Odrv4
    port map (
            O => \N__9442\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9439\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2111\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9430\
        );

    \I__2110\ : InMux
    port map (
            O => \N__9433\,
            I => \N__9427\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__9430\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__9427\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9422\,
            I => \N__9418\
        );

    \I__2106\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9415\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9418\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__9415\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__9410\,
            I => \N__9406\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9402\
        );

    \I__2101\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9399\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9405\,
            I => \N__9396\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9402\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__9399\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__9396\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2096\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9385\
        );

    \I__2095\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9382\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__9385\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__9382\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__9374\,
            I => \U409_TICK.TICK603_11\
        );

    \I__2090\ : InMux
    port map (
            O => \N__9371\,
            I => \N__9368\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9368\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2088\ : InMux
    port map (
            O => \N__9365\,
            I => \N__9361\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9358\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__9361\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2085\ : LocalMux
    port map (
            O => \N__9358\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2084\ : InMux
    port map (
            O => \N__9353\,
            I => \N__9350\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9350\,
            I => \U409_TICK.TICK503_11\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__9347\,
            I => \U409_TICK.TICK503_8_cascade_\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__9344\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__9341\,
            I => \N__9332\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__9340\,
            I => \N__9329\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9339\,
            I => \N__9319\
        );

    \I__2077\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9319\
        );

    \I__2076\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9319\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9336\,
            I => \N__9319\
        );

    \I__2074\ : InMux
    port map (
            O => \N__9335\,
            I => \N__9310\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9310\
        );

    \I__2072\ : InMux
    port map (
            O => \N__9329\,
            I => \N__9310\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9328\,
            I => \N__9310\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9319\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9310\,
            I => \U409_TICK.TICK503_9\
        );

    \I__2068\ : InMux
    port map (
            O => \N__9305\,
            I => \N__9299\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9304\,
            I => \N__9290\
        );

    \I__2066\ : InMux
    port map (
            O => \N__9303\,
            I => \N__9290\
        );

    \I__2065\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9290\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9299\,
            I => \N__9287\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9282\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9282\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9290\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2060\ : Odrv4
    port map (
            O => \N__9287\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9282\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2058\ : CascadeMux
    port map (
            O => \N__9275\,
            I => \N__9269\
        );

    \I__2057\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9263\
        );

    \I__2056\ : InMux
    port map (
            O => \N__9273\,
            I => \N__9256\
        );

    \I__2055\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9256\
        );

    \I__2054\ : InMux
    port map (
            O => \N__9269\,
            I => \N__9256\
        );

    \I__2053\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9253\
        );

    \I__2052\ : InMux
    port map (
            O => \N__9267\,
            I => \N__9248\
        );

    \I__2051\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9248\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__9263\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__9256\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9253\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__9248\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9227\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9227\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9227\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9236\,
            I => \N__9220\
        );

    \I__2042\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9220\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9234\,
            I => \N__9220\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9227\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__9220\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2038\ : CascadeMux
    port map (
            O => \N__9215\,
            I => \N__9209\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__9214\,
            I => \N__9206\
        );

    \I__2036\ : InMux
    port map (
            O => \N__9213\,
            I => \N__9202\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__9212\,
            I => \N__9199\
        );

    \I__2034\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9191\
        );

    \I__2033\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9191\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9205\,
            I => \N__9191\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9202\,
            I => \N__9188\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9183\
        );

    \I__2029\ : InMux
    port map (
            O => \N__9198\,
            I => \N__9183\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9191\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2027\ : Odrv4
    port map (
            O => \N__9188\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__9183\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9176\,
            I => \N__9172\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__9175\,
            I => \N__9168\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9165\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9162\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9159\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__9165\,
            I => \N__9154\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__9162\,
            I => \N__9154\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9159\,
            I => \N__9151\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__2016\ : Span4Mux_v
    port map (
            O => \N__9151\,
            I => \N__9143\
        );

    \I__2015\ : Span4Mux_h
    port map (
            O => \N__9148\,
            I => \N__9143\
        );

    \I__2014\ : Sp12to4
    port map (
            O => \N__9143\,
            I => \N__9140\
        );

    \I__2013\ : Odrv12
    port map (
            O => \N__9140\,
            I => \ROMEN\
        );

    \I__2012\ : IoInMux
    port map (
            O => \N__9137\,
            I => \N__9134\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__9134\,
            I => \N__9130\
        );

    \I__2010\ : IoInMux
    port map (
            O => \N__9133\,
            I => \N__9127\
        );

    \I__2009\ : IoSpan4Mux
    port map (
            O => \N__9130\,
            I => \N__9122\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9122\
        );

    \I__2007\ : IoSpan4Mux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__2006\ : IoSpan4Mux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__2005\ : Span4Mux_s0_v
    port map (
            O => \N__9116\,
            I => \N__9113\
        );

    \I__2004\ : Span4Mux_v
    port map (
            O => \N__9113\,
            I => \N__9109\
        );

    \I__2003\ : InMux
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__2002\ : Span4Mux_v
    port map (
            O => \N__9109\,
            I => \N__9101\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__9106\,
            I => \N__9101\
        );

    \I__2000\ : Span4Mux_v
    port map (
            O => \N__9101\,
            I => \N__9097\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9100\,
            I => \N__9094\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__9097\,
            I => \N__9091\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9088\
        );

    \I__1996\ : Odrv4
    port map (
            O => \N__9091\,
            I => \TACK_EN\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__9088\,
            I => \TACK_EN\
        );

    \I__1994\ : IoInMux
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__1992\ : Span4Mux_s2_v
    port map (
            O => \N__9077\,
            I => \N__9074\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__9071\,
            I => \N__9068\
        );

    \I__1989\ : Sp12to4
    port map (
            O => \N__9068\,
            I => \N__9065\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__9065\,
            I => \TCIn_1_i\
        );

    \I__1987\ : IoInMux
    port map (
            O => \N__9062\,
            I => \N__9059\
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9056\
        );

    \I__1985\ : Span4Mux_s3_v
    port map (
            O => \N__9056\,
            I => \N__9053\
        );

    \I__1984\ : Span4Mux_v
    port map (
            O => \N__9053\,
            I => \N__9050\
        );

    \I__1983\ : Span4Mux_h
    port map (
            O => \N__9050\,
            I => \N__9047\
        );

    \I__1982\ : Span4Mux_h
    port map (
            O => \N__9047\,
            I => \N__9043\
        );

    \I__1981\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9040\
        );

    \I__1980\ : Odrv4
    port map (
            O => \N__9043\,
            I => \TICK50_c\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__9040\,
            I => \TICK50_c\
        );

    \I__1978\ : InMux
    port map (
            O => \N__9035\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__1977\ : InMux
    port map (
            O => \N__9032\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9029\,
            I => \N__9025\
        );

    \I__1975\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9022\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__9025\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__9022\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9017\,
            I => \N__9013\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__9013\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__9010\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__9005\,
            I => \N__9002\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9002\,
            I => \N__8999\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__8999\,
            I => \N__8995\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8992\
        );

    \I__1964\ : Odrv4
    port map (
            O => \N__8995\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__8992\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__8987\,
            I => \N__8982\
        );

    \I__1961\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8979\
        );

    \I__1960\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8976\
        );

    \I__1959\ : InMux
    port map (
            O => \N__8982\,
            I => \N__8973\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8979\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8976\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8973\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__1955\ : InMux
    port map (
            O => \N__8966\,
            I => \N__8962\
        );

    \I__1954\ : InMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8962\,
            I => \N__8956\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__8959\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1951\ : Odrv12
    port map (
            O => \N__8956\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__1950\ : InMux
    port map (
            O => \N__8951\,
            I => \N__8948\
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8944\
        );

    \I__1948\ : InMux
    port map (
            O => \N__8947\,
            I => \N__8941\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__8944\,
            I => \N__8937\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__8941\,
            I => \N__8934\
        );

    \I__1945\ : InMux
    port map (
            O => \N__8940\,
            I => \N__8931\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__8937\,
            I => \U409_TRANSFER_ACK.N_101\
        );

    \I__1943\ : Odrv4
    port map (
            O => \N__8934\,
            I => \U409_TRANSFER_ACK.N_101\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8931\,
            I => \U409_TRANSFER_ACK.N_101\
        );

    \I__1941\ : InMux
    port map (
            O => \N__8924\,
            I => \N__8921\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8921\,
            I => \U409_TRANSFER_ACK.N_19\
        );

    \I__1939\ : IoInMux
    port map (
            O => \N__8918\,
            I => \N__8915\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__8915\,
            I => \N__8912\
        );

    \I__1937\ : Span4Mux_s0_v
    port map (
            O => \N__8912\,
            I => \N__8909\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__8909\,
            I => \N__8906\
        );

    \I__1935\ : Span4Mux_v
    port map (
            O => \N__8906\,
            I => \N__8903\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__8903\,
            I => \N__8899\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__8899\,
            I => \N__8890\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8887\
        );

    \I__1929\ : Odrv4
    port map (
            O => \N__8890\,
            I => \CLK_CIA_c\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__8887\,
            I => \CLK_CIA_c\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8882\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__1926\ : InMux
    port map (
            O => \N__8879\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__1925\ : InMux
    port map (
            O => \N__8876\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__1924\ : InMux
    port map (
            O => \N__8873\,
            I => \bfn_15_8_0_\
        );

    \I__1923\ : InMux
    port map (
            O => \N__8870\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8867\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8864\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8861\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8858\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__8855\,
            I => \U409_TRANSFER_ACK.N_19_cascade_\
        );

    \I__1917\ : InMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__8849\,
            I => \U409_TRANSFER_ACK.N_23\
        );

    \I__1915\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8843\,
            I => \U409_TRANSFER_ACK.N_22\
        );

    \I__1913\ : IoInMux
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1911\ : Span4Mux_s3_v
    port map (
            O => \N__8834\,
            I => \N__8831\
        );

    \I__1910\ : Sp12to4
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1909\ : Span12Mux_h
    port map (
            O => \N__8828\,
            I => \N__8824\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__1907\ : Odrv12
    port map (
            O => \N__8824\,
            I => \ROMENn_c\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8821\,
            I => \ROMENn_c\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8816\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__1904\ : InMux
    port map (
            O => \N__8813\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__1903\ : InMux
    port map (
            O => \N__8810\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8807\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8804\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__1900\ : InMux
    port map (
            O => \N__8801\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__1899\ : InMux
    port map (
            O => \N__8798\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8787\
        );

    \I__1897\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8784\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8793\,
            I => \N__8781\
        );

    \I__1895\ : InMux
    port map (
            O => \N__8792\,
            I => \N__8778\
        );

    \I__1894\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8773\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8790\,
            I => \N__8773\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__8787\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8784\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__8781\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8778\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8773\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__8762\,
            I => \N__8757\
        );

    \I__1886\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8753\
        );

    \I__1885\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8750\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8747\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8744\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__8753\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__8750\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8747\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__8744\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__8735\,
            I => \N__8730\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__8734\,
            I => \N__8726\
        );

    \I__1876\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8723\
        );

    \I__1875\ : InMux
    port map (
            O => \N__8730\,
            I => \N__8720\
        );

    \I__1874\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8717\
        );

    \I__1873\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8714\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__8723\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8720\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__8717\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__8714\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__8705\,
            I => \N__8697\
        );

    \I__1867\ : InMux
    port map (
            O => \N__8704\,
            I => \N__8692\
        );

    \I__1866\ : InMux
    port map (
            O => \N__8703\,
            I => \N__8692\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8702\,
            I => \N__8687\
        );

    \I__1864\ : InMux
    port map (
            O => \N__8701\,
            I => \N__8687\
        );

    \I__1863\ : InMux
    port map (
            O => \N__8700\,
            I => \N__8682\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8682\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__8692\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8687\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__8682\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8668\
        );

    \I__1857\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8663\
        );

    \I__1856\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8663\
        );

    \I__1855\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8660\
        );

    \I__1854\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8657\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__8668\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__8663\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__8660\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__8657\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1849\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__8645\,
            I => \U409_CIA.CLK_CIA6_0\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__8642\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_\
        );

    \I__1846\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8629\
        );

    \I__1845\ : InMux
    port map (
            O => \N__8638\,
            I => \N__8629\
        );

    \I__1844\ : InMux
    port map (
            O => \N__8637\,
            I => \N__8626\
        );

    \I__1843\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8623\
        );

    \I__1842\ : InMux
    port map (
            O => \N__8635\,
            I => \N__8618\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8618\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8629\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__8626\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__8623\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8618\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1835\ : LocalMux
    port map (
            O => \N__8606\,
            I => \N__8602\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8605\,
            I => \N__8599\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__8602\,
            I => \CIA_SPACE\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__8599\,
            I => \CIA_SPACE\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__8594\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8585\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0\
        );

    \I__1827\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8579\,
            I => \N__8573\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8570\
        );

    \I__1824\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8566\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8563\
        );

    \I__1822\ : Span4Mux_h
    port map (
            O => \N__8573\,
            I => \N__8558\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8558\
        );

    \I__1820\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8555\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8550\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8563\,
            I => \N__8550\
        );

    \I__1817\ : Span4Mux_h
    port map (
            O => \N__8558\,
            I => \N__8545\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8545\
        );

    \I__1815\ : Span4Mux_v
    port map (
            O => \N__8550\,
            I => \N__8542\
        );

    \I__1814\ : Span4Mux_v
    port map (
            O => \N__8545\,
            I => \N__8539\
        );

    \I__1813\ : Sp12to4
    port map (
            O => \N__8542\,
            I => \N__8534\
        );

    \I__1812\ : Sp12to4
    port map (
            O => \N__8539\,
            I => \N__8534\
        );

    \I__1811\ : Span12Mux_h
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1810\ : Span12Mux_v
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__8528\,
            I => \TSn_c\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__8525\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8522\,
            I => \N__8519\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8512\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8518\,
            I => \N__8512\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8517\,
            I => \N__8509\
        );

    \I__1803\ : LocalMux
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1801\ : Span4Mux_v
    port map (
            O => \N__8506\,
            I => \N__8500\
        );

    \I__1800\ : Span12Mux_h
    port map (
            O => \N__8503\,
            I => \N__8495\
        );

    \I__1799\ : Sp12to4
    port map (
            O => \N__8500\,
            I => \N__8495\
        );

    \I__1798\ : Odrv12
    port map (
            O => \N__8495\,
            I => \A_c_12\
        );

    \I__1797\ : IoInMux
    port map (
            O => \N__8492\,
            I => \N__8489\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__1795\ : IoSpan4Mux
    port map (
            O => \N__8486\,
            I => \N__8483\
        );

    \I__1794\ : Span4Mux_s3_h
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__1792\ : Span12Mux_h
    port map (
            O => \N__8477\,
            I => \N__8474\
        );

    \I__1791\ : Odrv12
    port map (
            O => \N__8474\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1790\ : InMux
    port map (
            O => \N__8471\,
            I => \N__8468\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8468\,
            I => \CIA_ENABLE\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8462\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8462\,
            I => \N__8457\
        );

    \I__1786\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8452\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8460\,
            I => \N__8452\
        );

    \I__1784\ : Span12Mux_v
    port map (
            O => \N__8457\,
            I => \N__8449\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__8452\,
            I => \N__8446\
        );

    \I__1782\ : Span12Mux_h
    port map (
            O => \N__8449\,
            I => \N__8443\
        );

    \I__1781\ : Span12Mux_v
    port map (
            O => \N__8446\,
            I => \N__8440\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__8443\,
            I => \A_c_13\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__8440\,
            I => \A_c_13\
        );

    \I__1778\ : IoInMux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1776\ : Span4Mux_s2_h
    port map (
            O => \N__8429\,
            I => \N__8426\
        );

    \I__1775\ : Sp12to4
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__1774\ : Span12Mux_s10_v
    port map (
            O => \N__8423\,
            I => \N__8420\
        );

    \I__1773\ : Odrv12
    port map (
            O => \N__8420\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__8417\,
            I => \N__8414\
        );

    \I__1771\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8408\
        );

    \I__1770\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8405\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8402\
        );

    \I__1768\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8399\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__8408\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__8405\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__8402\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8399\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8390\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8387\,
            I => \N__8376\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8376\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8376\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8373\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8370\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8376\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8373\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__8370\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__8363\,
            I => \N__8360\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8357\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8357\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\
        );

    \I__1751\ : InMux
    port map (
            O => \N__8354\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__1750\ : InMux
    port map (
            O => \N__8351\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8348\,
            I => \N__8345\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8345\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__8342\,
            I => \U409_CIA.CLK_CIA6_3_cascade_\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8339\,
            I => \N__8336\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__8336\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_2_1\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8330\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__8330\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__8327\,
            I => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\
        );

    \I__1741\ : InMux
    port map (
            O => \N__8324\,
            I => \N__8318\
        );

    \I__1740\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8318\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8318\,
            I => \U409_CIA.CIA_CLK_COUNT11_3\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__8315\,
            I => \U409_CIA.CLK_CIA6_0_cascade_\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8312\,
            I => \N__8309\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8309\,
            I => \U409_CIA.CLK_CIA6_3\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__8306\,
            I => \U409_CIA.CLK_CIA6_cascade_\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8303\,
            I => \N__8300\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8300\,
            I => \U409_CIA.CLK_CIA_RNOZ0Z_1\
        );

    \I__1732\ : InMux
    port map (
            O => \N__8297\,
            I => \N__8294\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8294\,
            I => \N__8290\
        );

    \I__1730\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8287\
        );

    \I__1729\ : Span4Mux_h
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__8287\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__8284\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__1726\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8275\
        );

    \I__1725\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8272\
        );

    \I__1724\ : LocalMux
    port map (
            O => \N__8275\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8272\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8267\,
            I => \N__8263\
        );

    \I__1721\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8260\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8263\,
            I => \N__8257\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8254\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__8257\,
            I => \N__8251\
        );

    \I__1717\ : Span4Mux_v
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1715\ : Sp12to4
    port map (
            O => \N__8248\,
            I => \N__8242\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__8245\,
            I => \N__8239\
        );

    \I__1713\ : Span12Mux_h
    port map (
            O => \N__8242\,
            I => \N__8236\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8239\,
            I => \N__8233\
        );

    \I__1711\ : Odrv12
    port map (
            O => \N__8236\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\
        );

    \I__1710\ : Odrv4
    port map (
            O => \N__8233\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\
        );

    \I__1709\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8224\
        );

    \I__1708\ : InMux
    port map (
            O => \N__8227\,
            I => \N__8221\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__8224\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8221\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8208\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8208\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8203\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8203\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__8208\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8203\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1699\ : CascadeMux
    port map (
            O => \N__8198\,
            I => \N__8194\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8197\,
            I => \N__8189\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8194\,
            I => \N__8184\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8184\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8192\,
            I => \N__8181\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8189\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8184\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8174\,
            I => \N__8167\
        );

    \I__1690\ : InMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8172\,
            I => \N__8164\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__8167\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__8164\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1686\ : IoInMux
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__1684\ : IoSpan4Mux
    port map (
            O => \N__8153\,
            I => \N__8150\
        );

    \I__1683\ : Span4Mux_s3_v
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1682\ : Sp12to4
    port map (
            O => \N__8147\,
            I => \N__8144\
        );

    \I__1681\ : Span12Mux_v
    port map (
            O => \N__8144\,
            I => \N__8140\
        );

    \I__1680\ : InMux
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8140\,
            I => \TACK_OUT\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__8137\,
            I => \TACK_OUT\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8132\,
            I => \N__8126\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8123\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8130\,
            I => \N__8118\
        );

    \I__1674\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8118\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__8126\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__8123\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__8118\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\
        );

    \I__1670\ : InMux
    port map (
            O => \N__8111\,
            I => \N__8106\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8110\,
            I => \N__8101\
        );

    \I__1668\ : InMux
    port map (
            O => \N__8109\,
            I => \N__8101\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8106\,
            I => \U409_TRANSFER_ACK.N_62\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__8101\,
            I => \U409_TRANSFER_ACK.N_62\
        );

    \I__1665\ : SRMux
    port map (
            O => \N__8096\,
            I => \N__8093\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__8093\,
            I => \N__8088\
        );

    \I__1663\ : SRMux
    port map (
            O => \N__8092\,
            I => \N__8085\
        );

    \I__1662\ : SRMux
    port map (
            O => \N__8091\,
            I => \N__8081\
        );

    \I__1661\ : Span4Mux_v
    port map (
            O => \N__8088\,
            I => \N__8078\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8075\
        );

    \I__1659\ : SRMux
    port map (
            O => \N__8084\,
            I => \N__8072\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8081\,
            I => \N__8069\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__8078\,
            I => \N__8064\
        );

    \I__1656\ : Span4Mux_v
    port map (
            O => \N__8075\,
            I => \N__8064\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8061\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__8069\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__8064\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1652\ : Odrv4
    port map (
            O => \N__8061\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8054\,
            I => \N__8051\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8051\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__8045\,
            I => \N__8038\
        );

    \I__1647\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8035\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8028\
        );

    \I__1645\ : InMux
    port map (
            O => \N__8042\,
            I => \N__8028\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8041\,
            I => \N__8025\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__8038\,
            I => \N__8020\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8035\,
            I => \N__8020\
        );

    \I__1641\ : InMux
    port map (
            O => \N__8034\,
            I => \N__8015\
        );

    \I__1640\ : InMux
    port map (
            O => \N__8033\,
            I => \N__8015\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__8028\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__8025\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1637\ : Odrv4
    port map (
            O => \N__8020\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__8015\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\
        );

    \I__1635\ : InMux
    port map (
            O => \N__8006\,
            I => \N__8002\
        );

    \I__1634\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7997\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8002\,
            I => \N__7994\
        );

    \I__1632\ : InMux
    port map (
            O => \N__8001\,
            I => \N__7991\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8000\,
            I => \N__7988\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__7997\,
            I => \N__7980\
        );

    \I__1629\ : Span4Mux_v
    port map (
            O => \N__7994\,
            I => \N__7980\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__7991\,
            I => \N__7980\
        );

    \I__1627\ : InMux
    port map (
            O => \N__7988\,
            I => \N__7975\
        );

    \I__1626\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7975\
        );

    \I__1625\ : Odrv4
    port map (
            O => \N__7980\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7975\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__1622\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7964\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7964\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__1620\ : IoInMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7955\
        );

    \I__1618\ : Span12Mux_s2_v
    port map (
            O => \N__7955\,
            I => \N__7952\
        );

    \I__1617\ : Odrv12
    port map (
            O => \N__7952\,
            I => \RESETn_c_i\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__7949\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7943\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7943\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\
        );

    \I__1613\ : InMux
    port map (
            O => \N__7940\,
            I => \N__7937\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7937\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\
        );

    \I__1611\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7930\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7933\,
            I => \N__7926\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__7930\,
            I => \N__7923\
        );

    \I__1608\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7920\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__7926\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1606\ : Odrv4
    port map (
            O => \N__7923\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7920\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__7913\,
            I => \N__7910\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1601\ : Odrv4
    port map (
            O => \N__7904\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7901\,
            I => \N__7891\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7891\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7899\,
            I => \N__7891\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7898\,
            I => \N__7888\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__7891\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7888\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__7883\,
            I => \N__7878\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7882\,
            I => \N__7872\
        );

    \I__1592\ : InMux
    port map (
            O => \N__7881\,
            I => \N__7869\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7878\,
            I => \N__7866\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7861\
        );

    \I__1589\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7861\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7858\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7872\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__7869\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__7866\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7861\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7858\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\
        );

    \I__1582\ : InMux
    port map (
            O => \N__7847\,
            I => \N__7840\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7846\,
            I => \N__7837\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7845\,
            I => \N__7832\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7844\,
            I => \N__7832\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7829\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7840\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__7837\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__7832\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__7829\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__7820\,
            I => \N__7814\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7811\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7818\,
            I => \N__7806\
        );

    \I__1570\ : InMux
    port map (
            O => \N__7817\,
            I => \N__7806\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7814\,
            I => \N__7803\
        );

    \I__1568\ : InMux
    port map (
            O => \N__7811\,
            I => \N__7800\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__7806\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7803\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__7800\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7793\,
            I => \N__7782\
        );

    \I__1563\ : InMux
    port map (
            O => \N__7792\,
            I => \N__7782\
        );

    \I__1562\ : InMux
    port map (
            O => \N__7791\,
            I => \N__7782\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7790\,
            I => \N__7777\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7789\,
            I => \N__7777\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__7782\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7777\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__7772\,
            I => \N__7769\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7762\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7767\,
            I => \N__7759\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7762\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7759\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\
        );

    \I__1551\ : IoInMux
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7748\
        );

    \I__1549\ : Span4Mux_s2_v
    port map (
            O => \N__7748\,
            I => \N__7745\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__7745\,
            I => \N__7742\
        );

    \I__1547\ : Odrv4
    port map (
            O => \N__7742\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__7739\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\
        );

    \I__1545\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7732\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7729\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7732\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__7729\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7724\,
            I => \N__7721\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7721\,
            I => \N__7717\
        );

    \I__1539\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__1538\ : Odrv12
    port map (
            O => \N__7717\,
            I => \AC_TACK\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__7714\,
            I => \AC_TACK\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__7709\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__7706\,
            I => \N__7703\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7703\,
            I => \N__7700\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7700\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\
        );

    \I__1532\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7691\
        );

    \I__1530\ : Span12Mux_h
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__1529\ : Span12Mux_v
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1528\ : Odrv12
    port map (
            O => \N__7685\,
            I => \CPUCONFn_c\
        );

    \I__1527\ : InMux
    port map (
            O => \N__7682\,
            I => \N__7679\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__7679\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__1525\ : InMux
    port map (
            O => \N__7676\,
            I => \N__7672\
        );

    \I__1524\ : InMux
    port map (
            O => \N__7675\,
            I => \N__7669\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7672\,
            I => \U409_AUTOCONFIG.STATE4\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7669\,
            I => \U409_AUTOCONFIG.STATE4\
        );

    \I__1521\ : InMux
    port map (
            O => \N__7664\,
            I => \N__7661\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__7661\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7655\,
            I => \N__7647\
        );

    \I__1517\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7642\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7642\
        );

    \I__1515\ : InMux
    port map (
            O => \N__7652\,
            I => \N__7639\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7651\,
            I => \N__7634\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7650\,
            I => \N__7634\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__7647\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7642\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7639\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__7634\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__7625\,
            I => \N__7617\
        );

    \I__1507\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7614\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__7623\,
            I => \N__7608\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__7622\,
            I => \N__7605\
        );

    \I__1504\ : InMux
    port map (
            O => \N__7621\,
            I => \N__7601\
        );

    \I__1503\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7598\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7617\,
            I => \N__7595\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__7614\,
            I => \N__7592\
        );

    \I__1500\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7589\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7612\,
            I => \N__7586\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7611\,
            I => \N__7579\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7579\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7605\,
            I => \N__7579\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__7604\,
            I => \N__7576\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7601\,
            I => \N__7569\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7569\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7595\,
            I => \N__7566\
        );

    \I__1491\ : Span4Mux_v
    port map (
            O => \N__7592\,
            I => \N__7561\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__7589\,
            I => \N__7561\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7558\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7579\,
            I => \N__7555\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7550\
        );

    \I__1486\ : InMux
    port map (
            O => \N__7575\,
            I => \N__7550\
        );

    \I__1485\ : InMux
    port map (
            O => \N__7574\,
            I => \N__7547\
        );

    \I__1484\ : Span4Mux_v
    port map (
            O => \N__7569\,
            I => \N__7542\
        );

    \I__1483\ : Span4Mux_v
    port map (
            O => \N__7566\,
            I => \N__7542\
        );

    \I__1482\ : Span4Mux_v
    port map (
            O => \N__7561\,
            I => \N__7539\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7558\,
            I => \N__7532\
        );

    \I__1480\ : Sp12to4
    port map (
            O => \N__7555\,
            I => \N__7532\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__7550\,
            I => \N__7532\
        );

    \I__1478\ : LocalMux
    port map (
            O => \N__7547\,
            I => \N__7525\
        );

    \I__1477\ : Sp12to4
    port map (
            O => \N__7542\,
            I => \N__7525\
        );

    \I__1476\ : Sp12to4
    port map (
            O => \N__7539\,
            I => \N__7525\
        );

    \I__1475\ : Span12Mux_h
    port map (
            O => \N__7532\,
            I => \N__7522\
        );

    \I__1474\ : Span12Mux_h
    port map (
            O => \N__7525\,
            I => \N__7519\
        );

    \I__1473\ : Span12Mux_v
    port map (
            O => \N__7522\,
            I => \N__7516\
        );

    \I__1472\ : Span12Mux_v
    port map (
            O => \N__7519\,
            I => \N__7513\
        );

    \I__1471\ : Odrv12
    port map (
            O => \N__7516\,
            I => \RnW_c\
        );

    \I__1470\ : Odrv12
    port map (
            O => \N__7513\,
            I => \RnW_c\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7508\,
            I => \N__7505\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7505\,
            I => \N__7497\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7504\,
            I => \N__7492\
        );

    \I__1466\ : InMux
    port map (
            O => \N__7503\,
            I => \N__7492\
        );

    \I__1465\ : InMux
    port map (
            O => \N__7502\,
            I => \N__7489\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7501\,
            I => \N__7486\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7500\,
            I => \N__7483\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__7497\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__7492\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__7489\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7486\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__7483\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1457\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__7469\,
            I => \N__7465\
        );

    \I__1455\ : InMux
    port map (
            O => \N__7468\,
            I => \N__7462\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__7465\,
            I => \N__7458\
        );

    \I__1453\ : LocalMux
    port map (
            O => \N__7462\,
            I => \N__7455\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7461\,
            I => \N__7452\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__7458\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__7455\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__7452\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7445\,
            I => \N__7441\
        );

    \I__1447\ : InMux
    port map (
            O => \N__7444\,
            I => \N__7438\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7441\,
            I => \N__7433\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7438\,
            I => \N__7433\
        );

    \I__1444\ : Span4Mux_v
    port map (
            O => \N__7433\,
            I => \N__7430\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__7430\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7424\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7424\,
            I => \N__7421\
        );

    \I__1440\ : Sp12to4
    port map (
            O => \N__7421\,
            I => \N__7418\
        );

    \I__1439\ : Span12Mux_v
    port map (
            O => \N__7418\,
            I => \N__7415\
        );

    \I__1438\ : Span12Mux_h
    port map (
            O => \N__7415\,
            I => \N__7412\
        );

    \I__1437\ : Odrv12
    port map (
            O => \N__7412\,
            I => \TACKn_in\
        );

    \I__1436\ : InMux
    port map (
            O => \N__7409\,
            I => \N__7406\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__7406\,
            I => \U409_TRANSFER_ACK.N_53\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__7403\,
            I => \U409_TRANSFER_ACK.N_53_cascade_\
        );

    \I__1433\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7397\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7397\,
            I => \N__7394\
        );

    \I__1431\ : Span4Mux_v
    port map (
            O => \N__7394\,
            I => \N__7390\
        );

    \I__1430\ : InMux
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__7390\,
            I => \ATA_SPACE\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__7387\,
            I => \ATA_SPACE\
        );

    \I__1427\ : IoInMux
    port map (
            O => \N__7382\,
            I => \N__7379\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__7379\,
            I => \N__7376\
        );

    \I__1425\ : Span12Mux_s3_v
    port map (
            O => \N__7376\,
            I => \N__7373\
        );

    \I__1424\ : Span12Mux_v
    port map (
            O => \N__7373\,
            I => \N__7370\
        );

    \I__1423\ : Span12Mux_h
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1422\ : Odrv12
    port map (
            O => \N__7367\,
            I => \BUFENn_c\
        );

    \I__1421\ : InMux
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7353\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7348\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7348\
        );

    \I__1417\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7345\
        );

    \I__1416\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7342\
        );

    \I__1415\ : InMux
    port map (
            O => \N__7356\,
            I => \N__7339\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__7353\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__7348\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__7345\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__7342\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7339\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__1409\ : IoInMux
    port map (
            O => \N__7328\,
            I => \N__7325\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7325\,
            I => \N__7322\
        );

    \I__1407\ : Span4Mux_s3_v
    port map (
            O => \N__7322\,
            I => \N__7319\
        );

    \I__1406\ : Span4Mux_v
    port map (
            O => \N__7319\,
            I => \N__7316\
        );

    \I__1405\ : Sp12to4
    port map (
            O => \N__7316\,
            I => \N__7313\
        );

    \I__1404\ : Span12Mux_h
    port map (
            O => \N__7313\,
            I => \N__7309\
        );

    \I__1403\ : InMux
    port map (
            O => \N__7312\,
            I => \N__7306\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__7309\,
            I => \CONFIGENn_c\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7306\,
            I => \CONFIGENn_c\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7301\,
            I => \N__7298\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7298\,
            I => \N__7290\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7287\
        );

    \I__1397\ : InMux
    port map (
            O => \N__7296\,
            I => \N__7284\
        );

    \I__1396\ : InMux
    port map (
            O => \N__7295\,
            I => \N__7277\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7294\,
            I => \N__7277\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7293\,
            I => \N__7277\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__7290\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__7287\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7284\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7277\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1389\ : InMux
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__7265\,
            I => \N__7260\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__7264\,
            I => \N__7257\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__7263\,
            I => \N__7251\
        );

    \I__1385\ : Span4Mux_v
    port map (
            O => \N__7260\,
            I => \N__7245\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7242\
        );

    \I__1383\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7237\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7237\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7254\,
            I => \N__7234\
        );

    \I__1380\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7225\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7225\
        );

    \I__1378\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7225\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7225\
        );

    \I__1376\ : Odrv4
    port map (
            O => \N__7245\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__7242\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7237\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__7234\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__7225\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7210\
        );

    \I__1370\ : InMux
    port map (
            O => \N__7213\,
            I => \N__7207\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7210\,
            I => \N__7204\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7207\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__7204\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__1366\ : InMux
    port map (
            O => \N__7199\,
            I => \N__7195\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7198\,
            I => \N__7192\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7187\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__7192\,
            I => \N__7187\
        );

    \I__1362\ : Span12Mux_v
    port map (
            O => \N__7187\,
            I => \N__7184\
        );

    \I__1361\ : Odrv12
    port map (
            O => \N__7184\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_13\
        );

    \I__1360\ : InMux
    port map (
            O => \N__7181\,
            I => \N__7178\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__1358\ : Span4Mux_h
    port map (
            O => \N__7175\,
            I => \N__7170\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7167\
        );

    \I__1356\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7164\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__7170\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1354\ : LocalMux
    port map (
            O => \N__7167\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7164\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__7157\,
            I => \N__7153\
        );

    \I__1351\ : CascadeMux
    port map (
            O => \N__7156\,
            I => \N__7149\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7153\,
            I => \N__7146\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7152\,
            I => \N__7143\
        );

    \I__1348\ : InMux
    port map (
            O => \N__7149\,
            I => \N__7138\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7146\,
            I => \N__7135\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7143\,
            I => \N__7132\
        );

    \I__1345\ : InMux
    port map (
            O => \N__7142\,
            I => \N__7129\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7126\
        );

    \I__1343\ : LocalMux
    port map (
            O => \N__7138\,
            I => \N__7121\
        );

    \I__1342\ : Span4Mux_v
    port map (
            O => \N__7135\,
            I => \N__7112\
        );

    \I__1341\ : Span4Mux_v
    port map (
            O => \N__7132\,
            I => \N__7112\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__7129\,
            I => \N__7112\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7112\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7125\,
            I => \N__7109\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__7124\,
            I => \N__7106\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__7121\,
            I => \N__7099\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__7112\,
            I => \N__7096\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__7109\,
            I => \N__7093\
        );

    \I__1333\ : InMux
    port map (
            O => \N__7106\,
            I => \N__7084\
        );

    \I__1332\ : InMux
    port map (
            O => \N__7105\,
            I => \N__7084\
        );

    \I__1331\ : InMux
    port map (
            O => \N__7104\,
            I => \N__7084\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7084\
        );

    \I__1329\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7081\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__7099\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__7096\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__7093\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7084\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__7081\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1323\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7067\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__7067\,
            I => \N__7059\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7066\,
            I => \N__7055\
        );

    \I__1320\ : InMux
    port map (
            O => \N__7065\,
            I => \N__7050\
        );

    \I__1319\ : InMux
    port map (
            O => \N__7064\,
            I => \N__7050\
        );

    \I__1318\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7047\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7062\,
            I => \N__7044\
        );

    \I__1316\ : Span4Mux_h
    port map (
            O => \N__7059\,
            I => \N__7041\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7058\,
            I => \N__7038\
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__7055\,
            I => \CONFIGURED\
        );

    \I__1313\ : LocalMux
    port map (
            O => \N__7050\,
            I => \CONFIGURED\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7047\,
            I => \CONFIGURED\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__7044\,
            I => \CONFIGURED\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__7041\,
            I => \CONFIGURED\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7038\,
            I => \CONFIGURED\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__7025\,
            I => \N__7020\
        );

    \I__1307\ : InMux
    port map (
            O => \N__7024\,
            I => \N__7013\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7023\,
            I => \N__7013\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7020\,
            I => \N__7013\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__7009\
        );

    \I__1303\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7006\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__7009\,
            I => \N__7003\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__7003\,
            I => \U409_AUTOCONFIG.N_192\
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__7000\,
            I => \U409_AUTOCONFIG.N_192\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6992\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6992\,
            I => \N__6989\
        );

    \I__1296\ : Odrv4
    port map (
            O => \N__6989\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_1\
        );

    \I__1295\ : CEMux
    port map (
            O => \N__6986\,
            I => \N__6982\
        );

    \I__1294\ : CEMux
    port map (
            O => \N__6985\,
            I => \N__6979\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6982\,
            I => \N__6975\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__6979\,
            I => \N__6972\
        );

    \I__1291\ : CEMux
    port map (
            O => \N__6978\,
            I => \N__6969\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__6975\,
            I => \N__6966\
        );

    \I__1289\ : Span4Mux_v
    port map (
            O => \N__6972\,
            I => \N__6963\
        );

    \I__1288\ : LocalMux
    port map (
            O => \N__6969\,
            I => \N__6960\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6966\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__6963\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1285\ : Odrv4
    port map (
            O => \N__6960\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__1283\ : InMux
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6947\,
            I => \N__6944\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__6944\,
            I => \U409_AUTOCONFIG.N_184_0\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6941\,
            I => \N__6935\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6935\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6935\,
            I => \U409_AUTOCONFIG.N_167\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6926\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6931\,
            I => \N__6926\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6926\,
            I => \U409_AUTOCONFIG.N_213_i\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6919\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6922\,
            I => \N__6915\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__6919\,
            I => \N__6912\
        );

    \I__1271\ : InMux
    port map (
            O => \N__6918\,
            I => \N__6909\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6915\,
            I => \U409_AUTOCONFIG.N_182_0\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__6912\,
            I => \U409_AUTOCONFIG.N_182_0\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6909\,
            I => \U409_AUTOCONFIG.N_182_0\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6896\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6896\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6896\,
            I => \N__6892\
        );

    \I__1264\ : InMux
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1263\ : Odrv4
    port map (
            O => \N__6892\,
            I => \U409_AUTOCONFIG.N_223\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__6889\,
            I => \U409_AUTOCONFIG.N_223\
        );

    \I__1261\ : InMux
    port map (
            O => \N__6884\,
            I => \N__6881\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6881\,
            I => \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__6878\,
            I => \N__6875\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6870\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6867\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6873\,
            I => \N__6864\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6870\,
            I => \N__6859\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__6867\,
            I => \N__6859\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6864\,
            I => \N__6853\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__6859\,
            I => \N__6850\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6858\,
            I => \N__6847\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6857\,
            I => \N__6844\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__6856\,
            I => \N__6841\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__6853\,
            I => \N__6837\
        );

    \I__1247\ : Span4Mux_v
    port map (
            O => \N__6850\,
            I => \N__6834\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6847\,
            I => \N__6829\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__6844\,
            I => \N__6829\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6824\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6840\,
            I => \N__6824\
        );

    \I__1242\ : Sp12to4
    port map (
            O => \N__6837\,
            I => \N__6821\
        );

    \I__1241\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6818\
        );

    \I__1240\ : Span4Mux_v
    port map (
            O => \N__6829\,
            I => \N__6813\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6824\,
            I => \N__6813\
        );

    \I__1238\ : Span12Mux_h
    port map (
            O => \N__6821\,
            I => \N__6810\
        );

    \I__1237\ : Span4Mux_v
    port map (
            O => \N__6818\,
            I => \N__6807\
        );

    \I__1236\ : Sp12to4
    port map (
            O => \N__6813\,
            I => \N__6804\
        );

    \I__1235\ : Span12Mux_v
    port map (
            O => \N__6810\,
            I => \N__6801\
        );

    \I__1234\ : Sp12to4
    port map (
            O => \N__6807\,
            I => \N__6796\
        );

    \I__1233\ : Span12Mux_v
    port map (
            O => \N__6804\,
            I => \N__6796\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6801\,
            I => \A_c_3\
        );

    \I__1231\ : Odrv12
    port map (
            O => \N__6796\,
            I => \A_c_3\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6788\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__6788\,
            I => \N__6785\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__6785\,
            I => \U409_AUTOCONFIG.N_190\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6773\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6770\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6765\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6779\,
            I => \N__6755\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6755\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6777\,
            I => \N__6750\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6776\,
            I => \N__6750\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6773\,
            I => \N__6745\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__6770\,
            I => \N__6745\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6740\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6740\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6737\
        );

    \I__1215\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6732\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6763\,
            I => \N__6732\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6729\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6724\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6724\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6715\
        );

    \I__1209\ : LocalMux
    port map (
            O => \N__6750\,
            I => \N__6715\
        );

    \I__1208\ : Span4Mux_h
    port map (
            O => \N__6745\,
            I => \N__6715\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6715\
        );

    \I__1206\ : Span4Mux_v
    port map (
            O => \N__6737\,
            I => \N__6712\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__6732\,
            I => \N__6707\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__6729\,
            I => \N__6707\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6724\,
            I => \N__6704\
        );

    \I__1202\ : Span4Mux_v
    port map (
            O => \N__6715\,
            I => \N__6701\
        );

    \I__1201\ : Span4Mux_v
    port map (
            O => \N__6712\,
            I => \N__6694\
        );

    \I__1200\ : Span4Mux_v
    port map (
            O => \N__6707\,
            I => \N__6694\
        );

    \I__1199\ : Span4Mux_v
    port map (
            O => \N__6704\,
            I => \N__6694\
        );

    \I__1198\ : Sp12to4
    port map (
            O => \N__6701\,
            I => \N__6689\
        );

    \I__1197\ : Sp12to4
    port map (
            O => \N__6694\,
            I => \N__6689\
        );

    \I__1196\ : Odrv12
    port map (
            O => \N__6689\,
            I => \A_c_4\
        );

    \I__1195\ : InMux
    port map (
            O => \N__6686\,
            I => \N__6680\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6680\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6668\
        );

    \I__1192\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6665\
        );

    \I__1191\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6662\
        );

    \I__1190\ : InMux
    port map (
            O => \N__6677\,
            I => \N__6657\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6657\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6675\,
            I => \N__6652\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6674\,
            I => \N__6652\
        );

    \I__1186\ : InMux
    port map (
            O => \N__6673\,
            I => \N__6647\
        );

    \I__1185\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6647\
        );

    \I__1184\ : InMux
    port map (
            O => \N__6671\,
            I => \N__6644\
        );

    \I__1183\ : Span4Mux_v
    port map (
            O => \N__6668\,
            I => \N__6631\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__6665\,
            I => \N__6631\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6662\,
            I => \N__6631\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__6657\,
            I => \N__6631\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6631\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6647\,
            I => \N__6626\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6644\,
            I => \N__6626\
        );

    \I__1176\ : InMux
    port map (
            O => \N__6643\,
            I => \N__6623\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6642\,
            I => \N__6620\
        );

    \I__1174\ : Span4Mux_v
    port map (
            O => \N__6631\,
            I => \N__6617\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6626\,
            I => \N__6614\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__6623\,
            I => \N__6609\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__6620\,
            I => \N__6609\
        );

    \I__1170\ : Sp12to4
    port map (
            O => \N__6617\,
            I => \N__6604\
        );

    \I__1169\ : Sp12to4
    port map (
            O => \N__6614\,
            I => \N__6604\
        );

    \I__1168\ : Span12Mux_h
    port map (
            O => \N__6609\,
            I => \N__6601\
        );

    \I__1167\ : Span12Mux_h
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__1166\ : Span12Mux_v
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__1165\ : Span12Mux_v
    port map (
            O => \N__6598\,
            I => \N__6592\
        );

    \I__1164\ : Odrv12
    port map (
            O => \N__6595\,
            I => \A_c_1\
        );

    \I__1163\ : Odrv12
    port map (
            O => \N__6592\,
            I => \A_c_1\
        );

    \I__1162\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6579\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6571\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6585\,
            I => \N__6571\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6584\,
            I => \N__6566\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6566\
        );

    \I__1157\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6563\
        );

    \I__1156\ : InMux
    port map (
            O => \N__6579\,
            I => \N__6559\
        );

    \I__1155\ : InMux
    port map (
            O => \N__6578\,
            I => \N__6556\
        );

    \I__1154\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6551\
        );

    \I__1153\ : InMux
    port map (
            O => \N__6576\,
            I => \N__6551\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__6571\,
            I => \N__6546\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__6566\,
            I => \N__6546\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6563\,
            I => \N__6543\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__6562\,
            I => \N__6540\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6533\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6556\,
            I => \N__6533\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__6551\,
            I => \N__6533\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__6546\,
            I => \N__6526\
        );

    \I__1144\ : Span4Mux_v
    port map (
            O => \N__6543\,
            I => \N__6523\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6520\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__6533\,
            I => \N__6517\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6532\,
            I => \N__6512\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6531\,
            I => \N__6512\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6507\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6507\
        );

    \I__1137\ : Sp12to4
    port map (
            O => \N__6526\,
            I => \N__6494\
        );

    \I__1136\ : Sp12to4
    port map (
            O => \N__6523\,
            I => \N__6494\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6520\,
            I => \N__6494\
        );

    \I__1134\ : Sp12to4
    port map (
            O => \N__6517\,
            I => \N__6494\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__6512\,
            I => \N__6494\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__6507\,
            I => \N__6494\
        );

    \I__1131\ : Span12Mux_h
    port map (
            O => \N__6494\,
            I => \N__6491\
        );

    \I__1130\ : Span12Mux_v
    port map (
            O => \N__6491\,
            I => \N__6488\
        );

    \I__1129\ : Odrv12
    port map (
            O => \N__6488\,
            I => \A_c_2\
        );

    \I__1128\ : InMux
    port map (
            O => \N__6485\,
            I => \N__6479\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6484\,
            I => \N__6476\
        );

    \I__1126\ : CascadeMux
    port map (
            O => \N__6483\,
            I => \N__6473\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__6482\,
            I => \N__6470\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6465\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6462\
        );

    \I__1122\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6457\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6470\,
            I => \N__6457\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__6469\,
            I => \N__6452\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6449\
        );

    \I__1118\ : Span4Mux_v
    port map (
            O => \N__6465\,
            I => \N__6442\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__6462\,
            I => \N__6442\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6457\,
            I => \N__6442\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6439\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6434\
        );

    \I__1113\ : InMux
    port map (
            O => \N__6452\,
            I => \N__6434\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6449\,
            I => \U409_AUTOCONFIG.N_198\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__6442\,
            I => \U409_AUTOCONFIG.N_198\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6439\,
            I => \U409_AUTOCONFIG.N_198\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__6434\,
            I => \U409_AUTOCONFIG.N_198\
        );

    \I__1108\ : InMux
    port map (
            O => \N__6425\,
            I => \N__6419\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6419\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1105\ : Odrv4
    port map (
            O => \N__6416\,
            I => \U409_AUTOCONFIG.N_222\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6413\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_\
        );

    \I__1103\ : IoInMux
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1101\ : IoSpan4Mux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1100\ : Sp12to4
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1099\ : Span12Mux_s7_v
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1098\ : Odrv12
    port map (
            O => \N__6395\,
            I => \D_OUT_0\
        );

    \I__1097\ : InMux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1095\ : Odrv12
    port map (
            O => \N__6386\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__1094\ : InMux
    port map (
            O => \N__6383\,
            I => \N__6380\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__6380\,
            I => \N__6377\
        );

    \I__1092\ : Odrv4
    port map (
            O => \N__6377\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6374\,
            I => \N__6365\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6365\
        );

    \I__1089\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6365\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6365\,
            I => \N__6361\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__6361\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6358\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1\
        );

    \I__1084\ : InMux
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1081\ : Sp12to4
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1080\ : Span12Mux_h
    port map (
            O => \N__6341\,
            I => \N__6338\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1078\ : Span12Mux_v
    port map (
            O => \N__6335\,
            I => \N__6332\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__6332\,
            I => \AUTOBOOT_c\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6326\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__6320\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_0\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6314\,
            I => \N__6311\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__6308\,
            I => \N__6304\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6301\
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__6304\,
            I => \U409_AUTOCONFIG.N_214_0\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6301\,
            I => \U409_AUTOCONFIG.N_214_0\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6290\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6290\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__6287\,
            I => \N__6282\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6279\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6285\,
            I => \N__6276\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__6282\,
            I => \U409_AUTOCONFIG.N_193_1\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6279\,
            I => \U409_AUTOCONFIG.N_193_1\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6276\,
            I => \U409_AUTOCONFIG.N_193_1\
        );

    \I__1056\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__6263\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__1053\ : InMux
    port map (
            O => \N__6260\,
            I => \N__6254\
        );

    \I__1052\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6254\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1050\ : Span4Mux_v
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1049\ : Odrv4
    port map (
            O => \N__6248\,
            I => \U409_AUTOCONFIG.N_159\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1047\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6239\,
            I => \N__6235\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__6238\,
            I => \N__6232\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__6235\,
            I => \N__6229\
        );

    \I__1043\ : InMux
    port map (
            O => \N__6232\,
            I => \N__6226\
        );

    \I__1042\ : Odrv4
    port map (
            O => \N__6229\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__6226\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6218\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1036\ : Odrv4
    port map (
            O => \N__6209\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__6200\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_2\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6197\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\
        );

    \I__1031\ : IoInMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__6191\,
            I => \N__6188\
        );

    \I__1029\ : Span12Mux_s8_v
    port map (
            O => \N__6188\,
            I => \N__6185\
        );

    \I__1028\ : Odrv12
    port map (
            O => \N__6185\,
            I => \D_OUT_2\
        );

    \I__1027\ : InMux
    port map (
            O => \N__6182\,
            I => \N__6174\
        );

    \I__1026\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6174\
        );

    \I__1025\ : CascadeMux
    port map (
            O => \N__6180\,
            I => \N__6171\
        );

    \I__1024\ : InMux
    port map (
            O => \N__6179\,
            I => \N__6167\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6164\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6171\,
            I => \N__6161\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6158\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6167\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10\
        );

    \I__1019\ : Odrv12
    port map (
            O => \N__6164\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6161\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__6158\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__6146\,
            I => \N__6143\
        );

    \I__1014\ : Span4Mux_h
    port map (
            O => \N__6143\,
            I => \N__6139\
        );

    \I__1013\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6136\
        );

    \I__1012\ : Span4Mux_v
    port map (
            O => \N__6139\,
            I => \N__6133\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__1010\ : Span4Mux_v
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1009\ : Span12Mux_h
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__1008\ : Odrv4
    port map (
            O => \N__6127\,
            I => \D_in_7\
        );

    \I__1007\ : Odrv12
    port map (
            O => \N__6124\,
            I => \D_in_7\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__6119\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_cascade_\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__6116\,
            I => \N__6113\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6110\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1002\ : Odrv12
    port map (
            O => \N__6107\,
            I => \U409_AUTOCONFIG.N_78\
        );

    \I__1001\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6100\
        );

    \I__1000\ : InMux
    port map (
            O => \N__6103\,
            I => \N__6091\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__6100\,
            I => \N__6088\
        );

    \I__998\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6085\
        );

    \I__997\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6082\
        );

    \I__996\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6075\
        );

    \I__995\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6075\
        );

    \I__994\ : InMux
    port map (
            O => \N__6095\,
            I => \N__6075\
        );

    \I__993\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6072\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6091\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__6088\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__6085\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__6082\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__6075\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__6072\,
            I => \U409_AUTOCONFIG.LIDE_BASE_10_2\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__6059\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_\
        );

    \I__985\ : IoInMux
    port map (
            O => \N__6056\,
            I => \N__6053\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__983\ : Span12Mux_s6_v
    port map (
            O => \N__6050\,
            I => \N__6047\
        );

    \I__982\ : Odrv12
    port map (
            O => \N__6047\,
            I => \D_OUT_1\
        );

    \I__981\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6041\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__979\ : InMux
    port map (
            O => \N__6038\,
            I => \N__6032\
        );

    \I__978\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6032\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__6032\,
            I => \U409_AUTOCONFIG.N_225\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6029\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_\
        );

    \I__975\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6023\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__6020\
        );

    \I__973\ : Odrv4
    port map (
            O => \N__6020\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3\
        );

    \I__972\ : InMux
    port map (
            O => \N__6017\,
            I => \N__6010\
        );

    \I__971\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6003\
        );

    \I__970\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6003\
        );

    \I__969\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6003\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__6013\,
            I => \N__5998\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__6010\,
            I => \N__5993\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6003\,
            I => \N__5993\
        );

    \I__965\ : InMux
    port map (
            O => \N__6002\,
            I => \N__5990\
        );

    \I__964\ : InMux
    port map (
            O => \N__6001\,
            I => \N__5985\
        );

    \I__963\ : InMux
    port map (
            O => \N__5998\,
            I => \N__5985\
        );

    \I__962\ : Span4Mux_v
    port map (
            O => \N__5993\,
            I => \N__5980\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5990\,
            I => \N__5980\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5985\,
            I => \N__5975\
        );

    \I__959\ : Sp12to4
    port map (
            O => \N__5980\,
            I => \N__5975\
        );

    \I__958\ : Odrv12
    port map (
            O => \N__5975\,
            I => \A_c_6\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__5972\,
            I => \N__5969\
        );

    \I__956\ : InMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5961\
        );

    \I__954\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5956\
        );

    \I__953\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5956\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__5961\,
            I => \N__5950\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__5956\,
            I => \N__5950\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__5955\,
            I => \N__5946\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__5950\,
            I => \N__5941\
        );

    \I__948\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5938\
        );

    \I__947\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5931\
        );

    \I__946\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5931\
        );

    \I__945\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5931\
        );

    \I__944\ : Sp12to4
    port map (
            O => \N__5941\,
            I => \N__5924\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5938\,
            I => \N__5924\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5931\,
            I => \N__5924\
        );

    \I__941\ : Span12Mux_h
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__5921\,
            I => \A_c_7\
        );

    \I__939\ : InMux
    port map (
            O => \N__5918\,
            I => \N__5914\
        );

    \I__938\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5911\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5911\,
            I => \U409_AUTOCONFIG.un1_A_13Z0Z_3\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__5908\,
            I => \U409_AUTOCONFIG.un1_A_13Z0Z_3\
        );

    \I__934\ : CascadeMux
    port map (
            O => \N__5903\,
            I => \U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_\
        );

    \I__933\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5897\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__5897\,
            I => \U409_AUTOCONFIG.N_70\
        );

    \I__931\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5890\
        );

    \I__930\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5887\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5890\,
            I => \LIDE_BASE_7\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__5887\,
            I => \LIDE_BASE_7\
        );

    \I__927\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5879\,
            I => \U409_AUTOCONFIG.N_74\
        );

    \I__925\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5872\
        );

    \I__924\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5868\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5872\,
            I => \N__5864\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__5871\,
            I => \N__5861\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5868\,
            I => \N__5858\
        );

    \I__920\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5855\
        );

    \I__919\ : Span4Mux_v
    port map (
            O => \N__5864\,
            I => \N__5850\
        );

    \I__918\ : InMux
    port map (
            O => \N__5861\,
            I => \N__5847\
        );

    \I__917\ : Span4Mux_v
    port map (
            O => \N__5858\,
            I => \N__5844\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__5855\,
            I => \N__5841\
        );

    \I__915\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5836\
        );

    \I__914\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5836\
        );

    \I__913\ : Sp12to4
    port map (
            O => \N__5850\,
            I => \N__5830\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5847\,
            I => \N__5830\
        );

    \I__911\ : Span4Mux_v
    port map (
            O => \N__5844\,
            I => \N__5827\
        );

    \I__910\ : Span4Mux_h
    port map (
            O => \N__5841\,
            I => \N__5822\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5836\,
            I => \N__5822\
        );

    \I__908\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5819\
        );

    \I__907\ : Span12Mux_h
    port map (
            O => \N__5830\,
            I => \N__5816\
        );

    \I__906\ : Span4Mux_v
    port map (
            O => \N__5827\,
            I => \N__5813\
        );

    \I__905\ : Sp12to4
    port map (
            O => \N__5822\,
            I => \N__5808\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5819\,
            I => \N__5808\
        );

    \I__903\ : Span12Mux_v
    port map (
            O => \N__5816\,
            I => \N__5805\
        );

    \I__902\ : Sp12to4
    port map (
            O => \N__5813\,
            I => \N__5800\
        );

    \I__901\ : Span12Mux_v
    port map (
            O => \N__5808\,
            I => \N__5800\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__5805\,
            I => \A_c_22\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__5800\,
            I => \A_c_22\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__5795\,
            I => \N__5789\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__5794\,
            I => \N__5786\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__5793\,
            I => \N__5783\
        );

    \I__895\ : InMux
    port map (
            O => \N__5792\,
            I => \N__5778\
        );

    \I__894\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5774\
        );

    \I__893\ : InMux
    port map (
            O => \N__5786\,
            I => \N__5767\
        );

    \I__892\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5764\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5761\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__5781\,
            I => \N__5758\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__5778\,
            I => \N__5755\
        );

    \I__888\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5752\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5774\,
            I => \N__5749\
        );

    \I__886\ : InMux
    port map (
            O => \N__5773\,
            I => \N__5746\
        );

    \I__885\ : InMux
    port map (
            O => \N__5772\,
            I => \N__5741\
        );

    \I__884\ : InMux
    port map (
            O => \N__5771\,
            I => \N__5741\
        );

    \I__883\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5737\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__5767\,
            I => \N__5732\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__5764\,
            I => \N__5732\
        );

    \I__880\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5729\
        );

    \I__879\ : InMux
    port map (
            O => \N__5758\,
            I => \N__5726\
        );

    \I__878\ : Span4Mux_h
    port map (
            O => \N__5755\,
            I => \N__5721\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5752\,
            I => \N__5721\
        );

    \I__876\ : Span4Mux_v
    port map (
            O => \N__5749\,
            I => \N__5714\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__5746\,
            I => \N__5714\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5714\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__5740\,
            I => \N__5711\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__5737\,
            I => \N__5702\
        );

    \I__871\ : Sp12to4
    port map (
            O => \N__5732\,
            I => \N__5702\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__5729\,
            I => \N__5702\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5726\,
            I => \N__5702\
        );

    \I__868\ : Span4Mux_v
    port map (
            O => \N__5721\,
            I => \N__5699\
        );

    \I__867\ : Span4Mux_v
    port map (
            O => \N__5714\,
            I => \N__5696\
        );

    \I__866\ : InMux
    port map (
            O => \N__5711\,
            I => \N__5693\
        );

    \I__865\ : Span12Mux_v
    port map (
            O => \N__5702\,
            I => \N__5684\
        );

    \I__864\ : Sp12to4
    port map (
            O => \N__5699\,
            I => \N__5684\
        );

    \I__863\ : Sp12to4
    port map (
            O => \N__5696\,
            I => \N__5684\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5684\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5684\,
            I => \A_c_21\
        );

    \I__860\ : CascadeMux
    port map (
            O => \N__5681\,
            I => \N__5678\
        );

    \I__859\ : InMux
    port map (
            O => \N__5678\,
            I => \N__5675\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5671\
        );

    \I__857\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__5671\,
            I => \LIDE_BASE_5\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__5668\,
            I => \LIDE_BASE_5\
        );

    \I__854\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5660\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5660\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\
        );

    \I__852\ : InMux
    port map (
            O => \N__5657\,
            I => \N__5654\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5654\,
            I => \N__5651\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__5651\,
            I => \U409_AUTOCONFIG.N_72\
        );

    \I__849\ : CascadeMux
    port map (
            O => \N__5648\,
            I => \N__5642\
        );

    \I__848\ : CascadeMux
    port map (
            O => \N__5647\,
            I => \N__5638\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__5646\,
            I => \N__5635\
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5645\,
            I => \N__5630\
        );

    \I__845\ : InMux
    port map (
            O => \N__5642\,
            I => \N__5623\
        );

    \I__844\ : InMux
    port map (
            O => \N__5641\,
            I => \N__5623\
        );

    \I__843\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5623\
        );

    \I__842\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5616\
        );

    \I__841\ : InMux
    port map (
            O => \N__5634\,
            I => \N__5616\
        );

    \I__840\ : InMux
    port map (
            O => \N__5633\,
            I => \N__5616\
        );

    \I__839\ : InMux
    port map (
            O => \N__5630\,
            I => \N__5613\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__5623\,
            I => \N__5610\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5616\,
            I => \U409_AUTOCONFIG.un1_STATE_6Z0Z_0\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__5613\,
            I => \U409_AUTOCONFIG.un1_STATE_6Z0Z_0\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__5610\,
            I => \U409_AUTOCONFIG.un1_STATE_6Z0Z_0\
        );

    \I__834\ : InMux
    port map (
            O => \N__5603\,
            I => \N__5597\
        );

    \I__833\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5597\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__5597\,
            I => \LIDE_BASE_6\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__830\ : InMux
    port map (
            O => \N__5591\,
            I => \N__5588\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__5588\,
            I => \N__5585\
        );

    \I__828\ : Odrv12
    port map (
            O => \N__5585\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_3\
        );

    \I__827\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__5576\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_0_2\
        );

    \I__824\ : InMux
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5570\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__822\ : InMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__820\ : Odrv12
    port map (
            O => \N__5561\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\
        );

    \I__819\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5551\
        );

    \I__818\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__817\ : InMux
    port map (
            O => \N__5556\,
            I => \N__5548\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__5551\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_5\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__5548\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_5\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5543\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_\
        );

    \I__813\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__5537\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1\
        );

    \I__811\ : IoInMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__809\ : IoSpan4Mux
    port map (
            O => \N__5528\,
            I => \N__5525\
        );

    \I__808\ : Span4Mux_s1_v
    port map (
            O => \N__5525\,
            I => \N__5522\
        );

    \I__807\ : Span4Mux_h
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__806\ : Sp12to4
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__805\ : Span12Mux_v
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__804\ : Odrv12
    port map (
            O => \N__5513\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__803\ : IoInMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5502\
        );

    \I__801\ : IoInMux
    port map (
            O => \N__5506\,
            I => \N__5499\
        );

    \I__800\ : IoInMux
    port map (
            O => \N__5505\,
            I => \N__5496\
        );

    \I__799\ : IoSpan4Mux
    port map (
            O => \N__5502\,
            I => \N__5493\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__5499\,
            I => \N__5488\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5496\,
            I => \N__5488\
        );

    \I__796\ : Span4Mux_s3_v
    port map (
            O => \N__5493\,
            I => \N__5482\
        );

    \I__795\ : Span4Mux_s3_v
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__794\ : IoInMux
    port map (
            O => \N__5487\,
            I => \N__5479\
        );

    \I__793\ : Span4Mux_v
    port map (
            O => \N__5482\,
            I => \N__5476\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__5476\,
            I => \D_1_i\
        );

    \I__790\ : Odrv12
    port map (
            O => \N__5473\,
            I => \D_1_i\
        );

    \I__789\ : InMux
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__787\ : Odrv12
    port map (
            O => \N__5462\,
            I => \D_in_4\
        );

    \I__786\ : InMux
    port map (
            O => \N__5459\,
            I => \N__5456\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5456\,
            I => \U409_AUTOCONFIG.N_76\
        );

    \I__784\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5447\
        );

    \I__783\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5447\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__781\ : Sp12to4
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__780\ : Span12Mux_v
    port map (
            O => \N__5441\,
            I => \N__5438\
        );

    \I__779\ : Odrv12
    port map (
            O => \N__5438\,
            I => \D_in_6\
        );

    \I__778\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5429\
        );

    \I__777\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5429\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__5426\,
            I => \N__5423\
        );

    \I__774\ : Span4Mux_v
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__5420\,
            I => \D_in_5\
        );

    \I__772\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__5414\,
            I => \U409_AUTOCONFIG.N_82\
        );

    \I__770\ : IoInMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__768\ : Span4Mux_s3_v
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__767\ : Span4Mux_v
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__5396\,
            I => \D_OUT_3\
        );

    \I__764\ : InMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5390\,
            I => \U409_AUTOCONFIG.N_80\
        );

    \I__762\ : CascadeMux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__761\ : InMux
    port map (
            O => \N__5384\,
            I => \N__5380\
        );

    \I__760\ : InMux
    port map (
            O => \N__5383\,
            I => \N__5377\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5380\,
            I => \LIDE_BASE_2\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__5377\,
            I => \LIDE_BASE_2\
        );

    \I__757\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5368\
        );

    \I__756\ : InMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5368\,
            I => \U409_ADDRESS_DECODE.N_34_1\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5365\,
            I => \U409_ADDRESS_DECODE.N_34_1\
        );

    \I__753\ : CascadeMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__752\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__5354\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0\
        );

    \I__750\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5347\
        );

    \I__749\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__5341\,
            I => \N__5333\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__5338\,
            I => \N__5333\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__5333\,
            I => \N_100\
        );

    \I__743\ : InMux
    port map (
            O => \N__5330\,
            I => \N__5327\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__5327\,
            I => \N__5323\
        );

    \I__741\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__740\ : Span12Mux_h
    port map (
            O => \N__5323\,
            I => \N__5314\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__5320\,
            I => \N__5314\
        );

    \I__738\ : InMux
    port map (
            O => \N__5319\,
            I => \N__5311\
        );

    \I__737\ : Odrv12
    port map (
            O => \N__5314\,
            I => \N_94\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__5311\,
            I => \N_94\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5306\,
            I => \U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_\
        );

    \I__734\ : IoInMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__732\ : Span4Mux_s3_v
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__730\ : Span4Mux_v
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__729\ : Span4Mux_v
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__728\ : Odrv4
    port map (
            O => \N__5285\,
            I => \PORTSIZE_0_i\
        );

    \I__727\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__5276\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0_0\
        );

    \I__724\ : InMux
    port map (
            O => \N__5273\,
            I => \N__5266\
        );

    \I__723\ : InMux
    port map (
            O => \N__5272\,
            I => \N__5257\
        );

    \I__722\ : InMux
    port map (
            O => \N__5271\,
            I => \N__5257\
        );

    \I__721\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5257\
        );

    \I__720\ : InMux
    port map (
            O => \N__5269\,
            I => \N__5257\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__5266\,
            I => \N__5254\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__717\ : Span4Mux_h
    port map (
            O => \N__5254\,
            I => \N__5247\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__5251\,
            I => \N__5244\
        );

    \I__715\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5241\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__5247\,
            I => \N__5238\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__5244\,
            I => \N__5233\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5241\,
            I => \N__5233\
        );

    \I__711\ : Sp12to4
    port map (
            O => \N__5238\,
            I => \N__5228\
        );

    \I__710\ : Span12Mux_h
    port map (
            O => \N__5233\,
            I => \N__5228\
        );

    \I__709\ : Odrv12
    port map (
            O => \N__5228\,
            I => \A_c_5\
        );

    \I__708\ : InMux
    port map (
            O => \N__5225\,
            I => \N__5221\
        );

    \I__707\ : InMux
    port map (
            O => \N__5224\,
            I => \N__5217\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5214\
        );

    \I__705\ : InMux
    port map (
            O => \N__5220\,
            I => \N__5211\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__5217\,
            I => \N__5206\
        );

    \I__703\ : Span4Mux_h
    port map (
            O => \N__5214\,
            I => \N__5200\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5200\
        );

    \I__701\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5197\
        );

    \I__700\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5194\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__5206\,
            I => \N__5191\
        );

    \I__698\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5188\
        );

    \I__697\ : Span4Mux_v
    port map (
            O => \N__5200\,
            I => \N__5179\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5179\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5194\,
            I => \N__5179\
        );

    \I__694\ : Span4Mux_v
    port map (
            O => \N__5191\,
            I => \N__5176\
        );

    \I__693\ : LocalMux
    port map (
            O => \N__5188\,
            I => \N__5173\
        );

    \I__692\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5170\
        );

    \I__691\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5167\
        );

    \I__690\ : Span4Mux_v
    port map (
            O => \N__5179\,
            I => \N__5164\
        );

    \I__689\ : Span4Mux_v
    port map (
            O => \N__5176\,
            I => \N__5157\
        );

    \I__688\ : Span4Mux_v
    port map (
            O => \N__5173\,
            I => \N__5157\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__5170\,
            I => \N__5157\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5167\,
            I => \N__5154\
        );

    \I__685\ : Sp12to4
    port map (
            O => \N__5164\,
            I => \N__5149\
        );

    \I__684\ : Sp12to4
    port map (
            O => \N__5157\,
            I => \N__5149\
        );

    \I__683\ : Span12Mux_v
    port map (
            O => \N__5154\,
            I => \N__5146\
        );

    \I__682\ : Odrv12
    port map (
            O => \N__5149\,
            I => \A_c_20\
        );

    \I__681\ : Odrv12
    port map (
            O => \N__5146\,
            I => \A_c_20\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__5141\,
            I => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_\
        );

    \I__679\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5132\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__5137\,
            I => \N__5129\
        );

    \I__677\ : CascadeMux
    port map (
            O => \N__5136\,
            I => \N__5124\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__5135\,
            I => \N__5121\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5132\,
            I => \N__5118\
        );

    \I__674\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5115\
        );

    \I__673\ : InMux
    port map (
            O => \N__5128\,
            I => \N__5110\
        );

    \I__672\ : InMux
    port map (
            O => \N__5127\,
            I => \N__5110\
        );

    \I__671\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5107\
        );

    \I__670\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5103\
        );

    \I__669\ : Span4Mux_v
    port map (
            O => \N__5118\,
            I => \N__5094\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5115\,
            I => \N__5094\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5094\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5107\,
            I => \N__5094\
        );

    \I__665\ : InMux
    port map (
            O => \N__5106\,
            I => \N__5091\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__5103\,
            I => \N__5088\
        );

    \I__663\ : Span4Mux_v
    port map (
            O => \N__5094\,
            I => \N__5083\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5091\,
            I => \N__5083\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__5088\,
            I => \N__5080\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__5083\,
            I => \N__5077\
        );

    \I__659\ : Sp12to4
    port map (
            O => \N__5080\,
            I => \N__5072\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__5077\,
            I => \N__5072\
        );

    \I__657\ : Odrv12
    port map (
            O => \N__5072\,
            I => \A_c_23\
        );

    \I__656\ : InMux
    port map (
            O => \N__5069\,
            I => \N__5063\
        );

    \I__655\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5063\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__5063\,
            I => \N__5058\
        );

    \I__653\ : InMux
    port map (
            O => \N__5062\,
            I => \N__5055\
        );

    \I__652\ : InMux
    port map (
            O => \N__5061\,
            I => \N__5052\
        );

    \I__651\ : Span4Mux_v
    port map (
            O => \N__5058\,
            I => \N__5047\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__5055\,
            I => \N__5047\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__5052\,
            I => \N__5044\
        );

    \I__648\ : Span4Mux_h
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__647\ : Span12Mux_v
    port map (
            O => \N__5044\,
            I => \N__5038\
        );

    \I__646\ : Odrv4
    port map (
            O => \N__5041\,
            I => \U409_ADDRESS_DECODE.N_92\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__5038\,
            I => \U409_ADDRESS_DECODE.N_92\
        );

    \I__644\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__5030\,
            I => \N__5026\
        );

    \I__642\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__5026\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_4\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__5023\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_4\
        );

    \I__639\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__5012\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE\
        );

    \I__636\ : InMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5006\,
            I => \U409_ADDRESS_DECODE.N_34\
        );

    \I__634\ : InMux
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5000\,
            I => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3\
        );

    \I__632\ : CascadeMux
    port map (
            O => \N__4997\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_cascade_\
        );

    \I__631\ : InMux
    port map (
            O => \N__4994\,
            I => \N__4991\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__4991\,
            I => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__4988\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__626\ : Odrv4
    port map (
            O => \N__4979\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4\
        );

    \I__625\ : CascadeMux
    port map (
            O => \N__4976\,
            I => \N__4972\
        );

    \I__624\ : InMux
    port map (
            O => \N__4975\,
            I => \N__4967\
        );

    \I__623\ : InMux
    port map (
            O => \N__4972\,
            I => \N__4967\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4967\,
            I => \U409_AUTOCONFIG.N_227_3\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__4964\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_\
        );

    \I__620\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4958\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4958\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__4955\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\
        );

    \I__617\ : InMux
    port map (
            O => \N__4952\,
            I => \N__4949\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4949\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__4946\,
            I => \ATA_SPACE_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__4943\,
            I => \N__4939\
        );

    \I__613\ : InMux
    port map (
            O => \N__4942\,
            I => \N__4936\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4939\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4936\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__610\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4924\
        );

    \I__608\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4921\
        );

    \I__607\ : Odrv12
    port map (
            O => \N__4924\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4921\,
            I => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\
        );

    \I__605\ : InMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4913\,
            I => \N__4908\
        );

    \I__603\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4905\
        );

    \I__602\ : InMux
    port map (
            O => \N__4911\,
            I => \N__4902\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__4908\,
            I => \N__4895\
        );

    \I__600\ : LocalMux
    port map (
            O => \N__4905\,
            I => \N__4895\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4902\,
            I => \N__4895\
        );

    \I__598\ : Span4Mux_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__596\ : Sp12to4
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__595\ : Span12Mux_h
    port map (
            O => \N__4886\,
            I => \N__4883\
        );

    \I__594\ : Odrv12
    port map (
            O => \N__4883\,
            I => \OVL_c\
        );

    \I__593\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4874\
        );

    \I__592\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4874\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4874\,
            I => \N__4869\
        );

    \I__590\ : InMux
    port map (
            O => \N__4873\,
            I => \N__4864\
        );

    \I__589\ : InMux
    port map (
            O => \N__4872\,
            I => \N__4864\
        );

    \I__588\ : Span4Mux_h
    port map (
            O => \N__4869\,
            I => \N__4858\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4864\,
            I => \N__4858\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__4863\,
            I => \N__4855\
        );

    \I__585\ : Span4Mux_v
    port map (
            O => \N__4858\,
            I => \N__4852\
        );

    \I__584\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4849\
        );

    \I__583\ : Sp12to4
    port map (
            O => \N__4852\,
            I => \N__4844\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4849\,
            I => \N__4844\
        );

    \I__581\ : Span12Mux_h
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__580\ : Span12Mux_v
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__579\ : Odrv12
    port map (
            O => \N__4838\,
            I => \A_c_19\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__4835\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_\
        );

    \I__577\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4829\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4824\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__4828\,
            I => \N__4821\
        );

    \I__574\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4818\
        );

    \I__573\ : Span4Mux_v
    port map (
            O => \N__4824\,
            I => \N__4813\
        );

    \I__572\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4810\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4818\,
            I => \N__4807\
        );

    \I__570\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4802\
        );

    \I__569\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4802\
        );

    \I__568\ : Sp12to4
    port map (
            O => \N__4813\,
            I => \N__4799\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4810\,
            I => \N__4796\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__4807\,
            I => \N__4791\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4802\,
            I => \N__4791\
        );

    \I__564\ : Span12Mux_s7_h
    port map (
            O => \N__4799\,
            I => \N__4786\
        );

    \I__563\ : Span12Mux_h
    port map (
            O => \N__4796\,
            I => \N__4786\
        );

    \I__562\ : Span4Mux_v
    port map (
            O => \N__4791\,
            I => \N__4783\
        );

    \I__561\ : Span12Mux_v
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__560\ : Sp12to4
    port map (
            O => \N__4783\,
            I => \N__4777\
        );

    \I__559\ : Odrv12
    port map (
            O => \N__4780\,
            I => \A_c_16\
        );

    \I__558\ : Odrv12
    port map (
            O => \N__4777\,
            I => \A_c_16\
        );

    \I__557\ : IoInMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4766\
        );

    \I__555\ : IoSpan4Mux
    port map (
            O => \N__4766\,
            I => \N__4763\
        );

    \I__554\ : Span4Mux_s2_v
    port map (
            O => \N__4763\,
            I => \N__4760\
        );

    \I__553\ : Span4Mux_v
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__552\ : Span4Mux_v
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__4754\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__550\ : InMux
    port map (
            O => \N__4751\,
            I => \N__4744\
        );

    \I__549\ : InMux
    port map (
            O => \N__4750\,
            I => \N__4744\
        );

    \I__548\ : InMux
    port map (
            O => \N__4749\,
            I => \N__4741\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4744\,
            I => \N__4735\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__4741\,
            I => \N__4732\
        );

    \I__545\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4729\
        );

    \I__544\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4726\
        );

    \I__543\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4723\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__4735\,
            I => \N__4720\
        );

    \I__541\ : Span4Mux_v
    port map (
            O => \N__4732\,
            I => \N__4717\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__4729\,
            I => \N__4714\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4726\,
            I => \N__4709\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__4723\,
            I => \N__4709\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__4720\,
            I => \N__4704\
        );

    \I__536\ : Sp12to4
    port map (
            O => \N__4717\,
            I => \N__4704\
        );

    \I__535\ : Span4Mux_v
    port map (
            O => \N__4714\,
            I => \N__4701\
        );

    \I__534\ : Span4Mux_v
    port map (
            O => \N__4709\,
            I => \N__4698\
        );

    \I__533\ : Span12Mux_s11_h
    port map (
            O => \N__4704\,
            I => \N__4695\
        );

    \I__532\ : Span4Mux_v
    port map (
            O => \N__4701\,
            I => \N__4692\
        );

    \I__531\ : Span4Mux_v
    port map (
            O => \N__4698\,
            I => \N__4689\
        );

    \I__530\ : Span12Mux_v
    port map (
            O => \N__4695\,
            I => \N__4682\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__4692\,
            I => \N__4682\
        );

    \I__528\ : Sp12to4
    port map (
            O => \N__4689\,
            I => \N__4682\
        );

    \I__527\ : Odrv12
    port map (
            O => \N__4682\,
            I => \A_c_18\
        );

    \I__526\ : InMux
    port map (
            O => \N__4679\,
            I => \N__4672\
        );

    \I__525\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__524\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4668\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4672\,
            I => \N__4665\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__4671\,
            I => \N__4662\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4668\,
            I => \N__4659\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__4665\,
            I => \N__4656\
        );

    \I__519\ : InMux
    port map (
            O => \N__4662\,
            I => \N__4653\
        );

    \I__518\ : Span12Mux_v
    port map (
            O => \N__4659\,
            I => \N__4650\
        );

    \I__517\ : Sp12to4
    port map (
            O => \N__4656\,
            I => \N__4645\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__4653\,
            I => \N__4645\
        );

    \I__515\ : Span12Mux_v
    port map (
            O => \N__4650\,
            I => \N__4642\
        );

    \I__514\ : Span12Mux_v
    port map (
            O => \N__4645\,
            I => \N__4639\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__4642\,
            I => \A_c_17\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__4639\,
            I => \A_c_17\
        );

    \I__511\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4628\
        );

    \I__510\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4628\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__4628\,
            I => \LIDE_BASE_1\
        );

    \I__508\ : InMux
    port map (
            O => \N__4625\,
            I => \N__4621\
        );

    \I__507\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4618\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4621\,
            I => \LIDE_BASE_4\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__4618\,
            I => \LIDE_BASE_4\
        );

    \I__504\ : InMux
    port map (
            O => \N__4613\,
            I => \N__4609\
        );

    \I__503\ : InMux
    port map (
            O => \N__4612\,
            I => \N__4606\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__4609\,
            I => \LIDE_BASE_3\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4606\,
            I => \LIDE_BASE_3\
        );

    \I__500\ : CascadeMux
    port map (
            O => \N__4601\,
            I => \N_89_cascade_\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4598\,
            I => \N_94_cascade_\
        );

    \I__498\ : InMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__496\ : Span4Mux_v
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__495\ : Odrv4
    port map (
            O => \N__4586\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1\
        );

    \I__494\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4580\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__492\ : Span4Mux_v
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__491\ : Span4Mux_h
    port map (
            O => \N__4574\,
            I => \N__4571\
        );

    \I__490\ : Sp12to4
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__489\ : Odrv12
    port map (
            O => \N__4568\,
            I => \TT_c_0\
        );

    \I__488\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__4559\,
            I => \N__4556\
        );

    \I__485\ : Span4Mux_h
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__483\ : Odrv12
    port map (
            O => \N__4550\,
            I => \TT_c_1\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__4547\,
            I => \N__4544\
        );

    \I__481\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4541\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__479\ : Odrv4
    port map (
            O => \N__4538\,
            I => \N_89\
        );

    \I__478\ : InMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__4532\,
            I => \N__4529\
        );

    \I__476\ : Odrv12
    port map (
            O => \N__4529\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__4526\,
            I => \N__4522\
        );

    \I__474\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4517\
        );

    \I__473\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4517\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__471\ : Span12Mux_v
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__470\ : Odrv12
    port map (
            O => \N__4511\,
            I => \A_c_15\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__4508\,
            I => \N__4505\
        );

    \I__468\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4499\
        );

    \I__467\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4499\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__465\ : Span4Mux_v
    port map (
            O => \N__4496\,
            I => \N__4493\
        );

    \I__464\ : Span4Mux_h
    port map (
            O => \N__4493\,
            I => \N__4490\
        );

    \I__463\ : Odrv4
    port map (
            O => \N__4490\,
            I => \A_c_25\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4487\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_\
        );

    \I__461\ : InMux
    port map (
            O => \N__4484\,
            I => \N__4478\
        );

    \I__460\ : InMux
    port map (
            O => \N__4483\,
            I => \N__4478\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__456\ : Sp12to4
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4466\,
            I => \A_c_24\
        );

    \I__454\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__4460\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\
        );

    \I__452\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__450\ : Span4Mux_v
    port map (
            O => \N__4451\,
            I => \N__4447\
        );

    \I__449\ : InMux
    port map (
            O => \N__4450\,
            I => \N__4444\
        );

    \I__448\ : Sp12to4
    port map (
            O => \N__4447\,
            I => \N__4439\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__4444\,
            I => \N__4439\
        );

    \I__446\ : Odrv12
    port map (
            O => \N__4439\,
            I => \A_c_27\
        );

    \I__445\ : InMux
    port map (
            O => \N__4436\,
            I => \N__4430\
        );

    \I__444\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4430\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__442\ : Span4Mux_v
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__441\ : Sp12to4
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__4421\,
            I => \A_c_30\
        );

    \I__439\ : CascadeMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__438\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4409\
        );

    \I__437\ : InMux
    port map (
            O => \N__4414\,
            I => \N__4409\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__435\ : Span4Mux_h
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__434\ : Span4Mux_v
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__433\ : Span4Mux_v
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__432\ : Odrv4
    port map (
            O => \N__4397\,
            I => \A_c_28\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__4394\,
            I => \N__4390\
        );

    \I__430\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4385\
        );

    \I__429\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4385\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__427\ : Sp12to4
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__426\ : Span12Mux_v
    port map (
            O => \N__4379\,
            I => \N__4376\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__4376\,
            I => \A_c_29\
        );

    \I__424\ : InMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__422\ : Span4Mux_v
    port map (
            O => \N__4367\,
            I => \N__4363\
        );

    \I__421\ : InMux
    port map (
            O => \N__4366\,
            I => \N__4360\
        );

    \I__420\ : Span4Mux_v
    port map (
            O => \N__4363\,
            I => \N__4357\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__4360\,
            I => \N__4354\
        );

    \I__418\ : Sp12to4
    port map (
            O => \N__4357\,
            I => \N__4351\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__4354\,
            I => \N__4348\
        );

    \I__416\ : Span12Mux_h
    port map (
            O => \N__4351\,
            I => \N__4343\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__4348\,
            I => \N__4343\
        );

    \I__414\ : Odrv12
    port map (
            O => \N__4343\,
            I => \A_c_31\
        );

    \I__413\ : InMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__4337\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__4334\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_\
        );

    \I__410\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__408\ : Odrv4
    port map (
            O => \N__4325\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10\
        );

    \I__407\ : IoInMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4319\,
            I => \N__4316\
        );

    \I__405\ : Span12Mux_s11_h
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__404\ : Span12Mux_h
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__403\ : Odrv12
    port map (
            O => \N__4310\,
            I => \N_61_i\
        );

    \I__402\ : IoInMux
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__401\ : LocalMux
    port map (
            O => \N__4304\,
            I => \N__4301\
        );

    \I__400\ : Span12Mux_s2_h
    port map (
            O => \N__4301\,
            I => \N__4298\
        );

    \I__399\ : Span12Mux_v
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__4295\,
            I => \SPIO_c\
        );

    \I__397\ : InMux
    port map (
            O => \N__4292\,
            I => \N__4286\
        );

    \I__396\ : InMux
    port map (
            O => \N__4291\,
            I => \N__4286\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__394\ : Span4Mux_v
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__393\ : Span4Mux_v
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__392\ : Sp12to4
    port map (
            O => \N__4277\,
            I => \N__4274\
        );

    \I__391\ : Odrv12
    port map (
            O => \N__4274\,
            I => \A_c_26\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__388\ : IoSpan4Mux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__387\ : Sp12to4
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__386\ : Span12Mux_s1_h
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__385\ : Span12Mux_v
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__384\ : Odrv12
    port map (
            O => \N__4253\,
            I => \PPIO_c\
        );

    \I__383\ : ClkMux
    port map (
            O => \N__4250\,
            I => \N__4211\
        );

    \I__382\ : ClkMux
    port map (
            O => \N__4249\,
            I => \N__4211\
        );

    \I__381\ : ClkMux
    port map (
            O => \N__4248\,
            I => \N__4211\
        );

    \I__380\ : ClkMux
    port map (
            O => \N__4247\,
            I => \N__4211\
        );

    \I__379\ : ClkMux
    port map (
            O => \N__4246\,
            I => \N__4211\
        );

    \I__378\ : ClkMux
    port map (
            O => \N__4245\,
            I => \N__4211\
        );

    \I__377\ : ClkMux
    port map (
            O => \N__4244\,
            I => \N__4211\
        );

    \I__376\ : ClkMux
    port map (
            O => \N__4243\,
            I => \N__4211\
        );

    \I__375\ : ClkMux
    port map (
            O => \N__4242\,
            I => \N__4211\
        );

    \I__374\ : ClkMux
    port map (
            O => \N__4241\,
            I => \N__4211\
        );

    \I__373\ : ClkMux
    port map (
            O => \N__4240\,
            I => \N__4211\
        );

    \I__372\ : ClkMux
    port map (
            O => \N__4239\,
            I => \N__4211\
        );

    \I__371\ : ClkMux
    port map (
            O => \N__4238\,
            I => \N__4211\
        );

    \I__370\ : GlobalMux
    port map (
            O => \N__4211\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__4250\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            I => \N__4249\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__4246\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4243\
        );

    \INVU409_TRANSFER_ACK.ROMENnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            I => \N__4248\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__4242\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__4240\
        );

    \INVU409_TRANSFER_ACK.TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            I => \N__4239\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__4238\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            I => \N__4245\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__4241\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__4247\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            I => \N__4244\
        );

    \INVU409_AUTOCONFIG.AC_TACKC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            I => \N__9889\
        );

    \INVU409_AUTOCONFIG.STATE_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_0C_net\,
            I => \N__9891\
        );

    \INVU409_AUTOCONFIG.CONFIGENnC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            I => \N__9898\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            I => \N__9896\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            I => \N__9895\
        );

    \INVU409_AUTOCONFIG.PR_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.PR_OUT_3C_net\,
            I => \N__9897\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_6C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_6C_net\,
            I => \N__9899\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\,
            I => \N__9904\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            I => \N__9905\
        );

    \IN_MUX_bfv_15_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_7_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_17_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_17_7_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7961\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_9_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4292\,
            in1 => \N__5351\,
            in2 => \N__4508\,
            in3 => \N__4484\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_3_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4291\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__4504\,
            in1 => \N__4463\,
            in2 => \N__4487\,
            in3 => \N__4483\,
            lcout => \U409_ADDRESS_DECODE.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a2_4_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4435\,
            in1 => \N__4366\,
            in2 => \N__4394\,
            in3 => \N__4414\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE_0_a2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_10_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4450\,
            in1 => \N__4436\,
            in2 => \N__4418\,
            in3 => \N__4393\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4749\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5186\,
            lcout => \N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_11_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4677\,
            in1 => \N__4535\,
            in2 => \N__5740\,
            in3 => \N__4373\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_tz_tz_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4595\,
            in1 => \N__4340\,
            in2 => \N__4334\,
            in3 => \N__4331\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_tz_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_61_i_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__4740\,
            in1 => \N__5326\,
            in2 => \N__5793\,
            in3 => \N__5220\,
            lcout => \N_61_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__6286\,
            in1 => \N__6781\,
            in2 => \N__6238\,
            in3 => \N__6582\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_0_0_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6468\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_0_1_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5792\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5210\,
            lcout => \U409_ADDRESS_DECODE.N_34_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_5_0_a3_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4879\,
            in1 => \N__4750\,
            in2 => \N__4828\,
            in3 => \N__4678\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4880\,
            in1 => \N__10412\,
            in2 => \N__5135\,
            in3 => \N__5875\,
            lcout => \N_89\,
            ltout => \N_89_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_i_a2_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__4679\,
            in1 => \_gnd_net_\,
            in2 => \N__4601\,
            in3 => \N__5062\,
            lcout => \N_94\,
            ltout => \N_94_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5209\,
            in1 => \N__5777\,
            in2 => \N__4598\,
            in3 => \N__4751\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14_8_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4583\,
            in1 => \N__4565\,
            in2 => \N__4547\,
            in3 => \N__4832\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_0_a3_0_14Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS0_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8460\,
            in1 => \N__4816\,
            in2 => \N__4526\,
            in3 => \N__8518\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS1_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__4817\,
            in1 => \N__4525\,
            in2 => \N__8522\,
            in3 => \N__8461\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_1_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__4738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5225\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_0_a2_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5770\,
            in1 => \N__5330\,
            in2 => \N__4835\,
            in3 => \N__4827\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__4931\,
            in1 => \N__4911\,
            in2 => \N__5794\,
            in3 => \N__5138\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__4739\,
            in1 => \N__5383\,
            in2 => \N__4671\,
            in3 => \N__4633\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_1_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000101010"
        )
    port map (
            in0 => \N__4634\,
            in1 => \N__6182\,
            in2 => \N__5647\,
            in3 => \N__5417\,
            lcout => \LIDE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__10130\
        );

    \U409_AUTOCONFIG.LIDE_BASE_3_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011111000000"
        )
    port map (
            in0 => \N__6181\,
            in1 => \N__5641\,
            in2 => \N__6116\,
            in3 => \N__4613\,
            lcout => \LIDE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__10130\
        );

    \U409_AUTOCONFIG.LIDE_BASE_4_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111000000"
        )
    port map (
            in0 => \N__6104\,
            in1 => \N__5459\,
            in2 => \N__5648\,
            in3 => \N__4625\,
            lcout => \LIDE_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__10130\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_4_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__5018\,
            in1 => \N__5893\,
            in2 => \N__5137\,
            in3 => \N__7058\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7214\,
            in1 => \N__5273\,
            in2 => \N__5972\,
            in3 => \N__5282\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__5224\,
            in1 => \N__4624\,
            in2 => \N__4863\,
            in3 => \N__4612\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4961\,
            in1 => \N__5663\,
            in2 => \N__4955\,
            in3 => \N__4952\,
            lcout => \ATA_SPACE\,
            ltout => \ATA_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__10393\,
            in1 => \N__7613\,
            in2 => \N__4946\,
            in3 => \N__4942\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9903\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__4927\,
            in1 => \N__5128\,
            in2 => \N__5782\,
            in3 => \N__4912\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__5867\,
            in1 => \N__5127\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7393\,
            in2 => \_gnd_net_\,
            in3 => \N__4943\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6456\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6643\,
            lcout => \U409_AUTOCONFIG.N_193_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000000"
        )
    port map (
            in0 => \N__5854\,
            in1 => \N__5069\,
            in2 => \N__10424\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.un1_RAMSPACEnZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_3_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__4873\,
            in1 => \N__4916\,
            in2 => \N__5781\,
            in3 => \N__5205\,
            lcout => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5853\,
            in1 => \N__5372\,
            in2 => \N__5136\,
            in3 => \N__4872\,
            lcout => \U409_ADDRESS_DECODE.N_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_14_2_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6578\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6780\,
            lcout => \U409_AUTOCONFIG.N_227_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.Z2_SPACE_0_a3_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__10420\,
            in1 => \N__5068\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE\,
            ltout => \U409_ADDRESS_DECODE.Z2_SPACE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__5009\,
            in1 => \N__5003\,
            in2 => \N__4997\,
            in3 => \N__4994\,
            lcout => \ROMEN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0_2_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__5945\,
            in1 => \N__6015\,
            in2 => \N__4976\,
            in3 => \N__5269\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_o3_2_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__6857\,
            in1 => \N__10394\,
            in2 => \N__4988\,
            in3 => \N__6672\,
            lcout => \U409_AUTOCONFIG.N_214_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4985\,
            in1 => \N__5272\,
            in2 => \N__5360\,
            in3 => \N__6762\,
            lcout => \U409_AUTOCONFIG.N_159\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_4_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__5944\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6014\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4\,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_2_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5271\,
            in1 => \N__4975\,
            in2 => \N__4964\,
            in3 => \N__6673\,
            lcout => \U409_AUTOCONFIG.N_192\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a2_1_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6858\,
            in1 => \N__5270\,
            in2 => \N__5955\,
            in3 => \N__6016\,
            lcout => \U409_AUTOCONFIG.N_198\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5371\,
            in1 => \N__5556\,
            in2 => \N__5871\,
            in3 => \N__5033\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6529\,
            in1 => \N__6840\,
            in2 => \_gnd_net_\,
            in3 => \N__6671\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PORTSIZE_1_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000111"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__5319\,
            in2 => \N__7156\,
            in3 => \N__5773\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.PORTSIZEZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PORTSIZE_0_i_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__10717\,
            in1 => \N__7461\,
            in2 => \N__5306\,
            in3 => \N__8605\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_STATE_6_0_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__6002\,
            in1 => \N__6761\,
            in2 => \N__6856\,
            in3 => \N__6530\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_3_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__6760\,
            in1 => \N__5250\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.un1_A_13Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_1_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5835\,
            in1 => \N__5187\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1\,
            ltout => \U409_ADDRESS_DECODE.un1_REGSPACEnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5771\,
            in1 => \N__5557\,
            in2 => \N__5141\,
            in3 => \N__5029\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_4_0_a3_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5106\,
            in1 => \N__5061\,
            in2 => \_gnd_net_\,
            in3 => \N__10413\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_4\,
            ltout => \U409_ADDRESS_DECODE.CIA_SPACE_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__5558\,
            in1 => \N__5772\,
            in2 => \N__5543\,
            in3 => \N__5540\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7624\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_4_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5468\,
            in1 => \N__7104\,
            in2 => \N__7622\,
            in3 => \N__6095\,
            lcout => \U409_AUTOCONFIG.N_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_6_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__6097\,
            in1 => \N__7611\,
            in2 => \N__7124\,
            in3 => \N__5453\,
            lcout => \U409_AUTOCONFIG.N_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_2_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6170\,
            in1 => \N__7125\,
            in2 => \N__7604\,
            in3 => \N__5452\,
            lcout => \U409_AUTOCONFIG.N_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_5_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5435\,
            in1 => \N__7105\,
            in2 => \N__7623\,
            in3 => \N__6096\,
            lcout => \U409_AUTOCONFIG.N_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_1_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5434\,
            in1 => \N__7575\,
            in2 => \N__6180\,
            in3 => \N__7103\,
            lcout => \U409_AUTOCONFIG.N_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__5567\,
            in1 => \N__7358\,
            in2 => \N__5594\,
            in3 => \N__7063\,
            lcout => \D_OUT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_2_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101011110000"
        )
    port map (
            in0 => \N__5393\,
            in1 => \N__6179\,
            in2 => \N__5387\,
            in3 => \N__5633\,
            lcout => \LIDE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\,
            ce => 'H',
            sr => \N__10129\
        );

    \U409_AUTOCONFIG.LIDE_BASE_7_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111000000"
        )
    port map (
            in0 => \N__6099\,
            in1 => \N__5900\,
            in2 => \N__5646\,
            in3 => \N__5894\,
            lcout => \LIDE_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\,
            ce => 'H',
            sr => \N__10129\
        );

    \U409_AUTOCONFIG.LIDE_BASE_5_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110011110000"
        )
    port map (
            in0 => \N__6098\,
            in1 => \N__5882\,
            in2 => \N__5681\,
            in3 => \N__5634\,
            lcout => \LIDE_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\,
            ce => 'H',
            sr => \N__10129\
        );

    \U409_AUTOCONFIG.CONFIGURED_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7181\,
            in1 => \N__7357\,
            in2 => \_gnd_net_\,
            in3 => \N__7062\,
            lcout => \CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_2C_net\,
            ce => 'H',
            sr => \N__10129\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__5876\,
            in1 => \N__5602\,
            in2 => \N__5795\,
            in3 => \N__5674\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_6_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111111000000"
        )
    port map (
            in0 => \N__6103\,
            in1 => \N__5657\,
            in2 => \N__5645\,
            in3 => \N__5603\,
            lcout => \LIDE_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_6C_net\,
            ce => 'H',
            sr => \N__10128\
        );

    \U409_AUTOCONFIG.PR_OUT_3_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__6026\,
            in1 => \N__10375\,
            in2 => \N__6587\,
            in3 => \N__6285\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.PR_OUT_3C_net\,
            ce => \N__6986\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_2_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10374\,
            in1 => \N__5582\,
            in2 => \_gnd_net_\,
            in3 => \N__7012\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.PR_OUT_3C_net\,
            ce => \N__6986\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__6364\,
            in1 => \N__6038\,
            in2 => \_gnd_net_\,
            in3 => \N__6922\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => \N__6978\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__6044\,
            in1 => \N__5573\,
            in2 => \_gnd_net_\,
            in3 => \N__7268\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6307\,
            in2 => \_gnd_net_\,
            in3 => \N__6037\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_3C_net\,
            ce => \N__6978\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_3_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__6577\,
            in1 => \N__6763\,
            in2 => \N__6469\,
            in3 => \N__6677\,
            lcout => \U409_AUTOCONFIG.N_225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_3_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6676\,
            in1 => \N__10377\,
            in2 => \N__6878\,
            in3 => \N__6576\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxa_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__6017\,
            in1 => \N__5949\,
            in2 => \N__6029\,
            in3 => \N__5917\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_0_sqmuxaZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6764\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6455\,
            lcout => \U409_AUTOCONFIG.PR_OUT_cnst_i_a4_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5964\,
            in1 => \N__6674\,
            in2 => \N__6013\,
            in3 => \N__6531\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_cnst_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_0_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__6675\,
            in1 => \N__6001\,
            in2 => \_gnd_net_\,
            in3 => \N__6874\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.un1_A_13Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5965\,
            in1 => \N__5918\,
            in2 => \N__5903\,
            in3 => \N__6532\,
            lcout => \U409_AUTOCONFIG.un1_AZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_7_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__6142\,
            in1 => \N__7141\,
            in2 => \N__7612\,
            in3 => \N__6094\,
            lcout => \U409_AUTOCONFIG.N_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7296\,
            in2 => \_gnd_net_\,
            in3 => \N__7254\,
            lcout => \U409_AUTOCONFIG.D_OUT_sm0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7250\,
            in1 => \N__6383\,
            in2 => \_gnd_net_\,
            in3 => \N__6269\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__6206\,
            in1 => \N__7360\,
            in2 => \N__6197\,
            in3 => \N__7065\,
            lcout => \D_OUT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6686\,
            in1 => \N__7294\,
            in2 => \_gnd_net_\,
            in3 => \N__7249\,
            lcout => \U409_AUTOCONFIG.LIDE_BASE_10\,
            ltout => \U409_AUTOCONFIG.LIDE_BASE_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_RNO_0_3_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6149\,
            in1 => \N__7142\,
            in2 => \N__6119\,
            in3 => \N__7621\,
            lcout => \U409_AUTOCONFIG.N_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNI0CVL_0_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6685\,
            in1 => \N__7293\,
            in2 => \_gnd_net_\,
            in3 => \N__7248\,
            lcout => \U409_AUTOCONFIG.LIDE_BASE_10_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIOO061_1_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__7295\,
            in1 => \N__6392\,
            in2 => \N__7263\,
            in3 => \N__6215\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_RNIOO061Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNID8KD2_1_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__6995\,
            in1 => \N__7359\,
            in2 => \N__6059\,
            in3 => \N__7064\,
            lcout => \D_OUT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIMM061_0_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101100"
        )
    port map (
            in0 => \N__6329\,
            in1 => \N__6221\,
            in2 => \N__7264\,
            in3 => \N__7301\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_RNIMM061Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIA5KD2_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__7364\,
            in1 => \N__6323\,
            in2 => \N__6413\,
            in3 => \N__7066\,
            lcout => \D_OUT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__6932\,
            in1 => \N__6373\,
            in2 => \N__10405\,
            in3 => \N__6296\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101110101010"
        )
    port map (
            in0 => \N__6374\,
            in1 => \N__6902\,
            in2 => \N__7025\,
            in3 => \N__6923\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110000010000"
        )
    port map (
            in0 => \N__6791\,
            in1 => \N__6372\,
            in2 => \N__6953\,
            in3 => \N__6353\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7023\,
            in1 => \N__6260\,
            in2 => \N__10403\,
            in3 => \N__6940\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__6901\,
            in1 => \N__6782\,
            in2 => \N__6317\,
            in3 => \N__6295\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000010"
        )
    port map (
            in0 => \N__10363\,
            in1 => \N__6259\,
            in2 => \N__6245\,
            in3 => \N__6931\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10364\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_1_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7024\,
            in1 => \N__6425\,
            in2 => \N__10404\,
            in3 => \N__6941\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_1C_net\,
            ce => \N__6985\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__7664\,
            in1 => \N__7502\,
            in2 => \N__10408\,
            in3 => \N__7675\,
            lcout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__6918\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6895\,
            lcout => \U409_AUTOCONFIG.N_184_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_a2_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6586\,
            in1 => \N__6779\,
            in2 => \_gnd_net_\,
            in3 => \N__6485\,
            lcout => \U409_AUTOCONFIG.N_167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_x3_0_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__6778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6585\,
            lcout => \U409_AUTOCONFIG.N_213_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_cnst_i_o3_3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001100"
        )
    port map (
            in0 => \N__6777\,
            in1 => \N__10376\,
            in2 => \N__6483\,
            in3 => \N__6584\,
            lcout => \U409_AUTOCONFIG.N_182_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_2_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__6776\,
            in1 => \N__6583\,
            in2 => \N__6482\,
            in3 => \N__6679\,
            lcout => \U409_AUTOCONFIG.N_223\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6769\,
            in1 => \N__6884\,
            in2 => \_gnd_net_\,
            in3 => \N__6873\,
            lcout => \U409_AUTOCONFIG.N_190\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_a3_1_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100000000"
        )
    port map (
            in0 => \N__6768\,
            in1 => \N__6678\,
            in2 => \N__6562\,
            in3 => \N__6484\,
            lcout => \U409_AUTOCONFIG.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LV_SPACE_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7444\,
            in1 => \N__7472\,
            in2 => \N__7157\,
            in3 => \N__7400\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__7356\,
            in1 => \N__7312\,
            in2 => \_gnd_net_\,
            in3 => \N__7173\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__10127\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7255\,
            in1 => \N__7174\,
            in2 => \_gnd_net_\,
            in3 => \N__7297\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__10127\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7199\,
            in1 => \N__7213\,
            in2 => \_gnd_net_\,
            in3 => \N__7256\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__10127\
        );

    \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7500\,
            in2 => \_gnd_net_\,
            in3 => \N__7650\,
            lcout => \U409_AUTOCONFIG.STATE_d_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__7651\,
            in1 => \N__7198\,
            in2 => \_gnd_net_\,
            in3 => \N__7501\,
            lcout => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__7503\,
            in1 => \N__7653\,
            in2 => \N__10406\,
            in3 => \N__7676\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000010100000"
        )
    port map (
            in0 => \N__7504\,
            in1 => \N__7620\,
            in2 => \N__10407\,
            in3 => \N__7654\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7152\,
            in1 => \N__8578\,
            in2 => \_gnd_net_\,
            in3 => \N__7070\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9890\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI04BC_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7682\,
            lcout => \U409_AUTOCONFIG.STATE4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__7574\,
            in1 => \N__7652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001000"
        )
    port map (
            in0 => \N__7720\,
            in1 => \N__7658\,
            in2 => \N__7625\,
            in3 => \N__7508\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__10124\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__7468\,
            in1 => \N__7445\,
            in2 => \N__10419\,
            in3 => \N__7427\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNO_0_5_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7881\,
            in2 => \_gnd_net_\,
            in3 => \N__7846\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_7_out\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110111011"
        )
    port map (
            in0 => \N__7736\,
            in1 => \N__7409\,
            in2 => \_gnd_net_\,
            in3 => \N__8110\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__8091\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_3_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__7876\,
            in1 => \N__8044\,
            in2 => \N__7706\,
            in3 => \N__7940\,
            lcout => \U409_TRANSFER_ACK.N_53\,
            ltout => \U409_TRANSFER_ACK.N_53_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQTP87_3_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111100001111"
        )
    port map (
            in0 => \N__9931\,
            in1 => \N__8569\,
            in2 => \N__7403\,
            in3 => \N__8109\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100001000"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__7934\,
            in2 => \N__7739\,
            in3 => \N__7847\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_ENC_net\,
            ce => 'H',
            sr => \N__8091\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__8048\,
            in1 => \N__8005\,
            in2 => \_gnd_net_\,
            in3 => \N__7790\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8084\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7929\,
            in1 => \N__7882\,
            in2 => \_gnd_net_\,
            in3 => \N__7789\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8084\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__8197\,
            in1 => \N__8216\,
            in2 => \N__10362\,
            in3 => \N__8172\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__10305\,
            in1 => \N__8192\,
            in2 => \_gnd_net_\,
            in3 => \N__8215\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_RNIGAOA_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8227\,
            in2 => \_gnd_net_\,
            in3 => \N__7735\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIBQIN_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__7724\,
            in1 => \N__8297\,
            in2 => \N__7709\,
            in3 => \N__8966\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__8034\,
            in1 => \N__8130\,
            in2 => \N__8000\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_0_7_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7898\,
            in1 => \N__7843\,
            in2 => \N__7819\,
            in3 => \N__7767\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_i_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI9U9R_2_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7987\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8129\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4\,
            ltout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER21_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIK98D3_0_3_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__8033\,
            in2 => \N__7949\,
            in3 => \N__7946\,
            lcout => \U409_TRANSFER_ACK.N_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__7817\,
            in1 => \N__7969\,
            in2 => \_gnd_net_\,
            in3 => \N__7792\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__8092\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI2DKM1_7_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7900\,
            in1 => \N__7844\,
            in2 => \N__7820\,
            in3 => \N__7768\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER23_i_0_o2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001101100"
        )
    port map (
            in0 => \N__7933\,
            in1 => \N__7901\,
            in2 => \N__7913\,
            in3 => \N__7791\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__8092\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNIQ4KM1_2_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7899\,
            in1 => \N__8131\,
            in2 => \N__7883\,
            in3 => \N__7845\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_ac0_9_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000001111000"
        )
    port map (
            in0 => \N__7818\,
            in1 => \N__7970\,
            in2 => \N__7772\,
            in3 => \N__7793\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6C_net\,
            ce => 'H',
            sr => \N__8092\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9933\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8582\,
            in1 => \N__8266\,
            in2 => \N__9935\,
            in3 => \N__8278\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000011110001"
        )
    port map (
            in0 => \N__8174\,
            in1 => \N__8193\,
            in2 => \N__9100\,
            in3 => \N__8213\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__10120\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__8947\,
            in1 => \N__8279\,
            in2 => \N__8267\,
            in3 => \N__8228\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__10120\
        );

    \U409_TRANSFER_ACK.TACK_OUT_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111011001010"
        )
    port map (
            in0 => \N__8214\,
            in1 => \N__8143\,
            in2 => \N__8198\,
            in3 => \N__8173\,
            lcout => \TACK_OUT\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_ENC_net\,
            ce => 'H',
            sr => \N__10120\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__8043\,
            in1 => \N__8132\,
            in2 => \_gnd_net_\,
            in3 => \N__8006\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__8096\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110000110011"
        )
    port map (
            in0 => \N__8576\,
            in1 => \N__8042\,
            in2 => \N__9934\,
            in3 => \N__8111\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__8096\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__8054\,
            in1 => \N__8041\,
            in2 => \_gnd_net_\,
            in3 => \N__8001\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10271\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001001011010"
        )
    port map (
            in0 => \N__8387\,
            in1 => \N__8333\,
            in2 => \N__8363\,
            in3 => \N__8324\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIMUMD1_7_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8756\,
            in1 => \N__8701\,
            in2 => \N__8734\,
            in3 => \N__8636\,
            lcout => \U409_CIA.CLK_CIA6_3\,
            ltout => \U409_CIA.CLK_CIA6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8672\,
            in1 => \N__8385\,
            in2 => \N__8342\,
            in3 => \N__8339\,
            lcout => \U409_CIA.CLK_CIA_RNOZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_2_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8790\,
            in2 => \_gnd_net_\,
            in3 => \N__8411\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIIQMD1_2_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__8386\,
            in1 => \N__8791\,
            in2 => \N__8417\,
            in3 => \N__8702\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_2_0\,
            ltout => \U409_CIA.CIA_CLK_COUNT11_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__8323\,
            in1 => \N__8795\,
            in2 => \N__8327\,
            in3 => \N__8348\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIQ2ND1_7_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8729\,
            in1 => \N__8637\,
            in2 => \N__8762\,
            in3 => \N__8674\,
            lcout => \U409_CIA.CIA_CLK_COUNT11_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNI9DRM_2_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8383\,
            in2 => \_gnd_net_\,
            in3 => \N__8413\,
            lcout => \U409_CIA.CLK_CIA6_0\,
            ltout => \U409_CIA.CLK_CIA6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8794\,
            in1 => \N__8673\,
            in2 => \N__8315\,
            in3 => \N__8312\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8895\,
            in2 => \N__8306\,
            in3 => \N__8303\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10910\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110100010"
        )
    port map (
            in0 => \N__8293\,
            in1 => \N__9213\,
            in2 => \N__8591\,
            in3 => \N__9305\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10121\
        );

    \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a4_1_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8577\,
            in2 => \_gnd_net_\,
            in3 => \N__9927\,
            lcout => \U409_TRANSFER_ACK.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_14_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10290\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10175\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8525\,
            in3 => \N__8517\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_14_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8471\,
            in2 => \_gnd_net_\,
            in3 => \N__8465\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8634\,
            in2 => \N__8705\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8412\,
            in2 => \_gnd_net_\,
            in3 => \N__8390\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__10911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_LUT4_0_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8384\,
            in2 => \_gnd_net_\,
            in3 => \N__8354\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8671\,
            in2 => \_gnd_net_\,
            in3 => \N__8351\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__10911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_LUT4_0_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8793\,
            in2 => \_gnd_net_\,
            in3 => \N__8804\,
            lcout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8761\,
            in2 => \_gnd_net_\,
            in3 => \N__8801\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__10911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8733\,
            in2 => \_gnd_net_\,
            in3 => \N__8798\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__8635\,
            in1 => \N__8700\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10911\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__8704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__8792\,
            in1 => \N__8760\,
            in2 => \N__8735\,
            in3 => \N__8703\,
            lcout => OPEN,
            ltout => \U409_CIA.un1_CIA_CLK_COUNT_3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_0_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000010000000"
        )
    port map (
            in0 => \N__8675\,
            in1 => \N__8648\,
            in2 => \N__8642\,
            in3 => \N__8638\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__8639\,
            in1 => \N__8609\,
            in2 => \N__8594\,
            in3 => \N__10164\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10909\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__9236\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9268\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER_5_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_1_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9298\,
            in1 => \N__9266\,
            in2 => \N__9212\,
            in3 => \N__9235\,
            lcout => \U409_TRANSFER_ACK.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI1MEE_1_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9234\,
            in1 => \N__9198\,
            in2 => \_gnd_net_\,
            in3 => \N__9297\,
            lcout => \U409_TRANSFER_ACK.N_19\,
            ltout => \U409_TRANSFER_ACK.N_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__8940\,
            in1 => \N__9171\,
            in2 => \N__8855\,
            in3 => \N__9267\,
            lcout => \U409_TRANSFER_ACK.N_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0000000011101110"
        )
    port map (
            in0 => \N__8827\,
            in1 => \N__8852\,
            in2 => \_gnd_net_\,
            in3 => \N__8846\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__10122\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9405\,
            in2 => \N__9487\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_15_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9421\,
            in2 => \_gnd_net_\,
            in3 => \N__8816\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__10786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9502\,
            in2 => \_gnd_net_\,
            in3 => \N__8813\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__10786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9364\,
            in2 => \_gnd_net_\,
            in3 => \N__8810\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9532\,
            in2 => \_gnd_net_\,
            in3 => \N__8807\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__10786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_15_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9445\,
            in2 => \_gnd_net_\,
            in3 => \N__8882\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_15_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8998\,
            in2 => \_gnd_net_\,
            in3 => \N__8879\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__10786\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9964\,
            in2 => \_gnd_net_\,
            in3 => \N__8876\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9679\,
            in2 => \_gnd_net_\,
            in3 => \N__8873\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9016\,
            in2 => \_gnd_net_\,
            in3 => \N__8870\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__10788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9517\,
            in2 => \_gnd_net_\,
            in3 => \N__8867\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__10788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9433\,
            in2 => \_gnd_net_\,
            in3 => \N__8864\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__10788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9028\,
            in2 => \_gnd_net_\,
            in3 => \N__8861\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__10788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9946\,
            in2 => \_gnd_net_\,
            in3 => \N__8858\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9805\,
            in2 => \_gnd_net_\,
            in3 => \N__9035\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9389\,
            in2 => \_gnd_net_\,
            in3 => \N__9032\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10788\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000001110000"
        )
    port map (
            in0 => \N__8986\,
            in1 => \N__9632\,
            in2 => \N__10402\,
            in3 => \N__9827\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9029\,
            in1 => \N__9017\,
            in2 => \N__9005\,
            in3 => \N__9806\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9965\,
            in1 => \N__9680\,
            in2 => \N__9452\,
            in3 => \N__9947\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000011001000"
        )
    port map (
            in0 => \N__8985\,
            in1 => \N__10361\,
            in2 => \N__9668\,
            in3 => \N__9818\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001001100"
        )
    port map (
            in0 => \N__9661\,
            in1 => \N__8965\,
            in2 => \N__8987\,
            in3 => \N__9836\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10125\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100000"
        )
    port map (
            in0 => \N__8951\,
            in1 => \N__9274\,
            in2 => \N__9175\,
            in3 => \N__8924\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10125\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8902\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__10125\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101110000"
        )
    port map (
            in0 => \N__9237\,
            in1 => \N__9205\,
            in2 => \N__9275\,
            in3 => \N__9302\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10123\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111110000000"
        )
    port map (
            in0 => \N__9304\,
            in1 => \N__9273\,
            in2 => \N__9215\,
            in3 => \N__9239\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10123\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011100001111000"
        )
    port map (
            in0 => \N__9303\,
            in1 => \N__9272\,
            in2 => \N__9214\,
            in3 => \N__9238\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__10123\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__9176\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9112\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9338\,
            in1 => \N__9588\,
            in2 => \N__10604\,
            in3 => \N__9625\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10065\,
            in1 => \_gnd_net_\,
            in2 => \N__10091\,
            in3 => \_gnd_net_\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_16_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9336\,
            in1 => \N__9586\,
            in2 => \N__10070\,
            in3 => \N__9623\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_16_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9585\,
            in1 => \N__9339\,
            in2 => \N__9626\,
            in3 => \N__9046\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9337\,
            in1 => \N__9587\,
            in2 => \N__9986\,
            in3 => \N__9624\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10787\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10043\,
            in1 => \N__10574\,
            in2 => \N__10090\,
            in3 => \N__10804\,
            lcout => \U409_TICK.TICK503_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_16_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10028\,
            in1 => \N__9998\,
            in2 => \_gnd_net_\,
            in3 => \N__10064\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_16_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9353\,
            in1 => \N__10499\,
            in2 => \N__9347\,
            in3 => \N__10535\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10013\,
            in1 => \N__10853\,
            in2 => \N__10592\,
            in3 => \N__10829\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9328\,
            in1 => \N__9590\,
            in2 => \N__9344\,
            in3 => \N__10508\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_16_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9589\,
            in1 => \N__9619\,
            in2 => \N__10841\,
            in3 => \N__9335\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_15_LC_16_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9617\,
            in1 => \N__9592\,
            in2 => \N__9340\,
            in3 => \N__10817\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_16_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9483\,
            in2 => \_gnd_net_\,
            in3 => \N__9409\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_16_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9618\,
            in1 => \N__9593\,
            in2 => \N__9341\,
            in3 => \N__10544\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_16_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10520\,
            in1 => \N__10556\,
            in2 => \N__10619\,
            in3 => \N__10484\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_16_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9616\,
            in1 => \N__9591\,
            in2 => \N__9560\,
            in3 => \N__10472\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10789\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__9714\,
            in1 => \N__9790\,
            in2 => \N__9767\,
            in3 => \N__9544\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__9533\,
            in1 => \N__9365\,
            in2 => \_gnd_net_\,
            in3 => \N__9482\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9377\,
            in1 => \N__9521\,
            in2 => \N__9506\,
            in3 => \N__9503\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__9488\,
            in1 => \N__9753\,
            in2 => \N__9491\,
            in3 => \N__9716\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9713\,
            in1 => \N__9789\,
            in2 => \N__9766\,
            in3 => \N__9458\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9434\,
            in1 => \N__9422\,
            in2 => \N__9410\,
            in3 => \N__9388\,
            lcout => \U409_TICK.TICK603_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9712\,
            in1 => \N__9788\,
            in2 => \N__9765\,
            in3 => \N__9371\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__9791\,
            in1 => \N__9715\,
            in2 => \N__9974\,
            in3 => \N__9763\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10791\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9792\,
            in1 => \N__9748\,
            in2 => \N__9724\,
            in3 => \N__9953\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__9932\,
            in1 => \N__10447\,
            in2 => \_gnd_net_\,
            in3 => \N__10462\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => \U409_TRANSFER_ACK.N_17_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101101011111"
        )
    port map (
            in0 => \N__9660\,
            in1 => \N__10434\,
            in2 => \N__9830\,
            in3 => \N__10145\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10448\,
            in2 => \_gnd_net_\,
            in3 => \N__10461\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => \U409_TRANSFER_ACK.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100100111"
        )
    port map (
            in0 => \N__9659\,
            in1 => \N__10435\,
            in2 => \N__9821\,
            in3 => \N__10146\,
            lcout => \U409_TRANSFER_ACK.N_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__9812\,
            in1 => \N__9720\,
            in2 => \N__9764\,
            in3 => \N__9794\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__9793\,
            in1 => \N__9749\,
            in2 => \N__9725\,
            in3 => \N__9686\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10793\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011100000100"
        )
    port map (
            in0 => \N__10147\,
            in1 => \N__9658\,
            in2 => \N__10439\,
            in3 => \N__9638\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10463\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__10126\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10148\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__10126\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10398\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10171\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__10126\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10083\,
            in2 => \N__10069\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10042\,
            in2 => \_gnd_net_\,
            in3 => \N__10031\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__10790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10027\,
            in2 => \_gnd_net_\,
            in3 => \N__10016\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__10790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10012\,
            in2 => \_gnd_net_\,
            in3 => \N__10001\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__10790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9997\,
            in2 => \_gnd_net_\,
            in3 => \N__9977\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10615\,
            in2 => \_gnd_net_\,
            in3 => \N__10595\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10588\,
            in2 => \_gnd_net_\,
            in3 => \N__10577\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__10790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10570\,
            in2 => \_gnd_net_\,
            in3 => \N__10559\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__10790\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10555\,
            in2 => \_gnd_net_\,
            in3 => \N__10538\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_7_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10534\,
            in2 => \_gnd_net_\,
            in3 => \N__10523\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__10792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10519\,
            in2 => \_gnd_net_\,
            in3 => \N__10502\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10498\,
            in2 => \_gnd_net_\,
            in3 => \N__10487\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__10792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10483\,
            in2 => \_gnd_net_\,
            in3 => \N__10466\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10852\,
            in2 => \_gnd_net_\,
            in3 => \N__10832\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10828\,
            in2 => \_gnd_net_\,
            in3 => \N__10811\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10805\,
            in2 => \_gnd_net_\,
            in3 => \N__10808\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__10792\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_0_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10727\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS1_LC_24_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10676\,
            lcout => \PCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS0_LC_24_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10672\,
            in2 => \_gnd_net_\,
            in3 => \N__10956\,
            lcout => \PCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS0_LC_24_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__10975\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10957\,
            lcout => \SCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS1_LC_24_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10958\,
            lcout => \SCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AGNUS_CLK_obuf_RNO_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10916\,
            in1 => \N__10889\,
            in2 => \_gnd_net_\,
            in3 => \N__10877\,
            lcout => \AGNUS_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

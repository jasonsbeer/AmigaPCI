-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 9 2025 18:43:01

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U111_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U111_TOP
entity U111_TOP is
port (
    D_UU_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_AMIGA : inout std_logic_vector(7 downto 0);
    D_UM_AMIGA : inout std_logic_vector(7 downto 0);
    D_LL_AMIGA : inout std_logic_vector(7 downto 0);
    D_LM_040 : inout std_logic_vector(7 downto 0);
    D_UM_040 : inout std_logic_vector(7 downto 0);
    D_LL_040 : inout std_logic_vector(7 downto 0);
    D_UU_040 : inout std_logic_vector(7 downto 0);
    A_AMIGA : out std_logic_vector(1 downto 0);
    A_040 : in std_logic_vector(1 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    TSn : out std_logic;
    RESETn : in std_logic;
    CLKRAMA : out std_logic;
    PORTSIZE : in std_logic;
    TEA_CPUn : out std_logic;
    LBENn : in std_logic;
    CLK40B : out std_logic;
    TBI_CPUn : out std_logic;
    TAn : inout std_logic;
    CPUBGn : out std_logic;
    BUFENn : out std_logic;
    RnW : in std_logic;
    CLK80_CPU : out std_logic;
    BUFDIR : out std_logic;
    TCI_CPUn : out std_logic;
    TS_CPUn : in std_logic;
    CLKRAMB : out std_logic;
    CLK40A : out std_logic;
    DMAn : out std_logic;
    CLK40C : out std_logic;
    CLK40_IN : in std_logic;
    TACKn : inout std_logic;
    BGn : in std_logic);
end U111_TOP;

-- Architecture of U111_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U111_TOP is

signal \N__8184\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8069\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8022\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__7997\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7968\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7932\ : std_logic;
signal \N__7925\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7898\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7896\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7887\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7871\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7860\ : std_logic;
signal \N__7853\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7842\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7815\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7790\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7752\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7727\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7716\ : std_logic;
signal \N__7709\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7664\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7628\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7599\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7581\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7572\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7563\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7536\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7527\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7502\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7465\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7446\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7376\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7374\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7365\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7356\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7347\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7281\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7272\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7263\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7257\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7230\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7190\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7170\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7112\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7095\ : std_logic;
signal \N__7092\ : std_logic;
signal \N__7089\ : std_logic;
signal \N__7086\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6837\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6758\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6681\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6630\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6612\ : std_logic;
signal \N__6609\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6459\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6449\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6339\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6198\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6144\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6122\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6072\ : std_logic;
signal \N__6069\ : std_logic;
signal \N__6066\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6009\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5819\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5766\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5664\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5621\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5603\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5586\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5382\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5352\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5313\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5190\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5162\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4987\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4872\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4861\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4858\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4855\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4819\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4816\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4614\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4455\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4422\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4410\ : std_logic;
signal \N__4407\ : std_logic;
signal \N__4404\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4339\ : std_logic;
signal \N__4336\ : std_logic;
signal \N__4333\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4318\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4312\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4231\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4197\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4140\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4134\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4125\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4096\ : std_logic;
signal \N__4093\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4078\ : std_logic;
signal \N__4075\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4057\ : std_logic;
signal \N__4056\ : std_logic;
signal \N__4053\ : std_logic;
signal \N__4050\ : std_logic;
signal \N__4047\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4041\ : std_logic;
signal \N__4038\ : std_logic;
signal \N__4035\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4026\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3988\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3894\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3873\ : std_logic;
signal \N__3870\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3859\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3853\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3829\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3808\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3802\ : std_logic;
signal \N__3799\ : std_logic;
signal \N__3796\ : std_logic;
signal \N__3793\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3730\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3724\ : std_logic;
signal \N__3721\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3717\ : std_logic;
signal \N__3714\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3702\ : std_logic;
signal \N__3699\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3646\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3640\ : std_logic;
signal \N__3637\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3633\ : std_logic;
signal \N__3630\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3583\ : std_logic;
signal \N__3580\ : std_logic;
signal \N__3577\ : std_logic;
signal \N__3574\ : std_logic;
signal \N__3571\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3526\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3442\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3426\ : std_logic;
signal \N__3423\ : std_logic;
signal \N__3420\ : std_logic;
signal \N__3417\ : std_logic;
signal \N__3414\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3396\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3316\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3310\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3283\ : std_logic;
signal \N__3280\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3223\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3205\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3190\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3174\ : std_logic;
signal \N__3171\ : std_logic;
signal \N__3168\ : std_logic;
signal \N__3165\ : std_logic;
signal \N__3162\ : std_logic;
signal \N__3159\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3150\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3142\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3136\ : std_logic;
signal \N__3133\ : std_logic;
signal \N__3130\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3121\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3111\ : std_logic;
signal \N__3108\ : std_logic;
signal \N__3105\ : std_logic;
signal \N__3102\ : std_logic;
signal \N__3099\ : std_logic;
signal \N__3096\ : std_logic;
signal \N__3093\ : std_logic;
signal \N__3088\ : std_logic;
signal \N__3085\ : std_logic;
signal \N__3082\ : std_logic;
signal \N__3079\ : std_logic;
signal \N__3076\ : std_logic;
signal \N__3073\ : std_logic;
signal \N__3070\ : std_logic;
signal \N__3067\ : std_logic;
signal \N__3064\ : std_logic;
signal \N__3061\ : std_logic;
signal \N__3058\ : std_logic;
signal \N__3055\ : std_logic;
signal \N__3052\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3043\ : std_logic;
signal \N__3040\ : std_logic;
signal \N__3037\ : std_logic;
signal \N__3034\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3028\ : std_logic;
signal \N__3025\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3010\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2983\ : std_logic;
signal \N__2980\ : std_logic;
signal \N__2979\ : std_logic;
signal \N__2976\ : std_logic;
signal \N__2973\ : std_logic;
signal \N__2970\ : std_logic;
signal \N__2967\ : std_logic;
signal \N__2964\ : std_logic;
signal \N__2961\ : std_logic;
signal \N__2958\ : std_logic;
signal \N__2955\ : std_logic;
signal \N__2952\ : std_logic;
signal \N__2949\ : std_logic;
signal \N__2946\ : std_logic;
signal \N__2943\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2935\ : std_logic;
signal \N__2932\ : std_logic;
signal \N__2929\ : std_logic;
signal \N__2926\ : std_logic;
signal \N__2923\ : std_logic;
signal \N__2920\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2914\ : std_logic;
signal \N__2911\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2859\ : std_logic;
signal \N__2856\ : std_logic;
signal \N__2853\ : std_logic;
signal \N__2850\ : std_logic;
signal \N__2847\ : std_logic;
signal \N__2842\ : std_logic;
signal \N__2839\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2830\ : std_logic;
signal \N__2827\ : std_logic;
signal \N__2824\ : std_logic;
signal \N__2821\ : std_logic;
signal \N__2818\ : std_logic;
signal \N__2815\ : std_logic;
signal \N__2814\ : std_logic;
signal \N__2811\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2767\ : std_logic;
signal \N__2764\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2758\ : std_logic;
signal \N__2755\ : std_logic;
signal \N__2752\ : std_logic;
signal \N__2749\ : std_logic;
signal \N__2746\ : std_logic;
signal \N__2745\ : std_logic;
signal \N__2742\ : std_logic;
signal \N__2739\ : std_logic;
signal \N__2736\ : std_logic;
signal \N__2733\ : std_logic;
signal \N__2730\ : std_logic;
signal \N__2727\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2718\ : std_logic;
signal \N__2715\ : std_logic;
signal \N__2712\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2701\ : std_logic;
signal \N__2698\ : std_logic;
signal \N__2695\ : std_logic;
signal \N__2692\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2686\ : std_logic;
signal \N__2683\ : std_logic;
signal \N__2680\ : std_logic;
signal \N__2677\ : std_logic;
signal \N__2674\ : std_logic;
signal \N__2671\ : std_logic;
signal \N__2668\ : std_logic;
signal \N__2665\ : std_logic;
signal \N__2662\ : std_logic;
signal \N__2659\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2653\ : std_logic;
signal \N__2650\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2644\ : std_logic;
signal \N__2641\ : std_logic;
signal \N__2638\ : std_logic;
signal \N__2635\ : std_logic;
signal \N__2632\ : std_logic;
signal \N__2629\ : std_logic;
signal \N__2626\ : std_logic;
signal \N__2623\ : std_logic;
signal \N__2620\ : std_logic;
signal \N__2617\ : std_logic;
signal \N__2614\ : std_logic;
signal \N__2611\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2605\ : std_logic;
signal \N__2602\ : std_logic;
signal \N__2599\ : std_logic;
signal \N__2596\ : std_logic;
signal \N__2593\ : std_logic;
signal \N__2590\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2574\ : std_logic;
signal \N__2573\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2569\ : std_logic;
signal \N__2566\ : std_logic;
signal \N__2563\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2559\ : std_logic;
signal \N__2558\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2546\ : std_logic;
signal \N__2543\ : std_logic;
signal \N__2542\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2531\ : std_logic;
signal \N__2530\ : std_logic;
signal \N__2529\ : std_logic;
signal \N__2526\ : std_logic;
signal \N__2523\ : std_logic;
signal \N__2520\ : std_logic;
signal \N__2517\ : std_logic;
signal \N__2514\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2512\ : std_logic;
signal \N__2511\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2509\ : std_logic;
signal \N__2508\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2496\ : std_logic;
signal \N__2493\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2489\ : std_logic;
signal \N__2488\ : std_logic;
signal \N__2485\ : std_logic;
signal \N__2482\ : std_logic;
signal \N__2479\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2475\ : std_logic;
signal \N__2474\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2472\ : std_logic;
signal \N__2469\ : std_logic;
signal \N__2468\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2460\ : std_logic;
signal \N__2457\ : std_logic;
signal \N__2454\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2452\ : std_logic;
signal \N__2451\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2449\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2437\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2431\ : std_logic;
signal \N__2428\ : std_logic;
signal \N__2425\ : std_logic;
signal \N__2422\ : std_logic;
signal \N__2419\ : std_logic;
signal \N__2412\ : std_logic;
signal \N__2409\ : std_logic;
signal \N__2406\ : std_logic;
signal \N__2403\ : std_logic;
signal \N__2400\ : std_logic;
signal \N__2397\ : std_logic;
signal \N__2396\ : std_logic;
signal \N__2395\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2366\ : std_logic;
signal \N__2363\ : std_logic;
signal \N__2360\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2340\ : std_logic;
signal \N__2337\ : std_logic;
signal \N__2334\ : std_logic;
signal \N__2331\ : std_logic;
signal \N__2326\ : std_logic;
signal \N__2323\ : std_logic;
signal \N__2320\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TAn_in\ : std_logic;
signal \A_040_c_1\ : std_logic;
signal \A_040_c_0\ : std_logic;
signal \A_AMIGA_c_0\ : std_logic;
signal \RnW_c_i\ : std_logic;
signal \D_LL_040_in_2\ : std_logic;
signal \D_UM_040_in_2\ : std_logic;
signal \un1_D_UM_040_2\ : std_logic;
signal \D_LM_AMIGA_in_5\ : std_logic;
signal \un1_D_LM_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_6\ : std_logic;
signal \un1_D_LM_AMIGA_6\ : std_logic;
signal \D_LL_040_in_3\ : std_logic;
signal \D_UM_040_in_3\ : std_logic;
signal \un1_D_UM_040_3\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \D_UU_040_in_6\ : std_logic;
signal \D_LM_040_in_6\ : std_logic;
signal \un1_D_UU_040_6\ : std_logic;
signal \D_UU_040_in_0\ : std_logic;
signal \D_LM_040_in_0\ : std_logic;
signal \un1_D_UU_040_0\ : std_logic;
signal \D_LM_AMIGA_in_3\ : std_logic;
signal \un1_D_LM_AMIGA_3\ : std_logic;
signal \D_LM_AMIGA_in_2\ : std_logic;
signal \un1_D_LM_AMIGA_2\ : std_logic;
signal \D_LL_040_in_7\ : std_logic;
signal \D_UM_040_in_7\ : std_logic;
signal \un1_D_UM_040_7\ : std_logic;
signal \D_LL_AMIGA_in_0\ : std_logic;
signal \un1_D_LL_AMIGA_0\ : std_logic;
signal \LBENn_c_i_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \INVU111_CYCLE_SM.TSnC_net\ : std_logic;
signal \D_LL_AMIGA_in_5\ : std_logic;
signal \un1_D_LL_AMIGA_5\ : std_logic;
signal \D_LM_AMIGA_in_4\ : std_logic;
signal \un1_D_LM_AMIGA_4\ : std_logic;
signal \D_UM_040_in_6\ : std_logic;
signal \D_LL_040_in_6\ : std_logic;
signal \un1_D_UM_040_6\ : std_logic;
signal \D_LL_040_in_1\ : std_logic;
signal \D_UM_040_in_1\ : std_logic;
signal \un1_D_UM_040_1\ : std_logic;
signal \LBENn_c_i\ : std_logic;
signal \D_LM_040_in_1\ : std_logic;
signal \D_UU_040_in_1\ : std_logic;
signal \un1_D_UU_040_1\ : std_logic;
signal \D_LM_040_in_4\ : std_logic;
signal \D_UU_040_in_4\ : std_logic;
signal \un1_D_UU_040_4\ : std_logic;
signal \D_UU_040_in_2\ : std_logic;
signal \D_LM_040_in_2\ : std_logic;
signal \un1_D_UU_040_2\ : std_logic;
signal \D_LL_AMIGA_in_2\ : std_logic;
signal \un1_D_LL_AMIGA_2\ : std_logic;
signal \D_LL_AMIGA_in_4\ : std_logic;
signal \un1_D_LL_AMIGA_4\ : std_logic;
signal \D_LL_AMIGA_in_6\ : std_logic;
signal \un1_D_LL_AMIGA_6\ : std_logic;
signal \D_LM_AMIGA_in_0\ : std_logic;
signal \un1_D_LM_AMIGA_0\ : std_logic;
signal \D_LL_AMIGA_in_7\ : std_logic;
signal \un1_D_LL_AMIGA_7\ : std_logic;
signal \D_LL_040_in_0\ : std_logic;
signal \D_UM_040_in_0\ : std_logic;
signal \un1_D_UM_040_0\ : std_logic;
signal \D_UM_040_in_4\ : std_logic;
signal \D_LL_040_in_4\ : std_logic;
signal \un1_D_UM_040_4\ : std_logic;
signal \D_LM_040_in_5\ : std_logic;
signal \D_UU_040_in_5\ : std_logic;
signal \un1_D_UU_040_5\ : std_logic;
signal \D_LM_040_in_7\ : std_logic;
signal \D_UU_040_in_7\ : std_logic;
signal \un1_D_UU_040_7\ : std_logic;
signal \D_LL_AMIGA_in_3\ : std_logic;
signal \un1_D_LL_AMIGA_3\ : std_logic;
signal \D_LL_AMIGA_in_1\ : std_logic;
signal \un1_D_LL_AMIGA_1\ : std_logic;
signal \A_AMIGA_c_1\ : std_logic;
signal \D_LM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.FLIP_cascade_\ : std_logic;
signal \un1_D_LM_AMIGA_1\ : std_logic;
signal \GB_BUFFER_CLK40_THRU_CO\ : std_logic;
signal \CLK80\ : std_logic;
signal \GB_BUFFER_CLK80_THRU_CO\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.A_OUTZ0\ : std_logic;
signal \U111_CYCLE_SM.N_75_0_cascade_\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\ : std_logic;
signal \U111_CYCLE_SM.TS_ENZ0\ : std_logic;
signal \U111_CYCLE_SM.un3_LW_CYCLE_START\ : std_logic;
signal \INVU111_CYCLE_SM.TA_ENC_net\ : std_logic;
signal \U111_CYCLE_SM.RESETn_c_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \PORTSIZE_c\ : std_logic;
signal \U111_CYCLE_SM.LW_TRANS_0\ : std_logic;
signal \D_LM_AMIGA_in_7\ : std_logic;
signal \un1_D_LM_AMIGA_7\ : std_logic;
signal \D_LL_040_in_5\ : std_logic;
signal \D_UM_040_in_5\ : std_logic;
signal \un1_D_UM_040_5\ : std_logic;
signal \D_UU_040_in_3\ : std_logic;
signal \U111_CYCLE_SM.FLIP\ : std_logic;
signal \D_LM_040_in_3\ : std_logic;
signal \un1_D_UU_040_3\ : std_logic;
signal \U111_CYCLE_SM_TBI_CPUn_0_i\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_5\ : std_logic;
signal \BGn_c\ : std_logic;
signal \CPU_READ_EN_i\ : std_logic;
signal \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\ : std_logic;
signal \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_STARTZ0\ : std_logic;
signal \U111_CYCLE_SM.N_97_cascade_\ : std_logic;
signal \INVU111_CYCLE_SM.LW_CYCLEC_net\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLE_0\ : std_logic;
signal \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\ : std_logic;
signal \D_UU_AMIGA_in_1\ : std_logic;
signal \un1_D_UU_AMIGA_1\ : std_logic;
signal \U111_CYCLE_SM.TA_ENZ0\ : std_logic;
signal \LBENn_c\ : std_logic;
signal \TAn_1_i\ : std_logic;
signal \D_UM_AMIGA_in_1\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\ : std_logic;
signal \un1_D_UM_AMIGA_1\ : std_logic;
signal \TS_CPUn_c\ : std_logic;
signal \CLK40\ : std_logic;
signal \U111_CYCLE_SM.TS_EN_2_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\ : std_logic;
signal \D_UU_AMIGA_in_7\ : std_logic;
signal \un1_D_UU_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\ : std_logic;
signal \D_UU_AMIGA_in_2\ : std_logic;
signal \un1_D_UU_AMIGA_2\ : std_logic;
signal \un1_D_UM_AMIGA_0\ : std_logic;
signal \un1_D_UM_AMIGA_2\ : std_logic;
signal \un1_D_UM_AMIGA_6\ : std_logic;
signal \D_UM_AMIGA_in_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\ : std_logic;
signal \D_UM_AMIGA_in_6\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\ : std_logic;
signal \D_UM_AMIGA_in_2\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\ : std_logic;
signal \D_UM_AMIGA_in_5\ : std_logic;
signal \un1_D_UM_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\ : std_logic;
signal \D_UU_AMIGA_in_3\ : std_logic;
signal \un1_D_UU_AMIGA_3\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\ : std_logic;
signal \D_UU_AMIGA_in_4\ : std_logic;
signal \un1_D_UU_AMIGA_4\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\ : std_logic;
signal \D_UU_AMIGA_in_6\ : std_logic;
signal \un1_D_UU_AMIGA_6\ : std_logic;
signal \D_UM_AMIGA_in_3\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\ : std_logic;
signal \un1_D_UM_AMIGA_3\ : std_logic;
signal \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\ : std_logic;
signal \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\ : std_logic;
signal \D_UM_AMIGA_in_7\ : std_logic;
signal \un1_D_UM_AMIGA_7\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\ : std_logic;
signal \D_UU_AMIGA_in_0\ : std_logic;
signal \un1_D_UU_AMIGA_0\ : std_logic;
signal \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\ : std_logic;
signal \D_UU_AMIGA_in_5\ : std_logic;
signal \un1_D_UU_AMIGA_5\ : std_logic;
signal \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\ : std_logic;
signal \D_UM_AMIGA_in_4\ : std_logic;
signal \U111_CYCLE_SM.LW_CYCLEZ0\ : std_logic;
signal \un1_D_UM_AMIGA_4\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \LBENn_wire\ : std_logic;
signal \CPUBGn_wire\ : std_logic;
signal \TEA_CPUn_wire\ : std_logic;
signal \A_040_wire\ : std_logic_vector(1 downto 0);
signal \A_AMIGA_wire\ : std_logic_vector(1 downto 0);
signal \CLK40B_wire\ : std_logic;
signal \BUFDIR_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \TS_CPUn_wire\ : std_logic;
signal \CLKRAMA_wire\ : std_logic;
signal \TCI_CPUn_wire\ : std_logic;
signal \CLKRAMB_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \DMAn_wire\ : std_logic;
signal \CLK80_CPU_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40C_wire\ : std_logic;
signal \BGn_wire\ : std_logic;
signal \TBI_CPUn_wire\ : std_logic;
signal \CLK40A_wire\ : std_logic;
signal \pll_pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \LBENn_wire\ <= LBENn;
    CPUBGn <= \CPUBGn_wire\;
    TEA_CPUn <= \TEA_CPUn_wire\;
    \A_040_wire\ <= A_040;
    A_AMIGA <= \A_AMIGA_wire\;
    CLK40B <= \CLK40B_wire\;
    BUFDIR <= \BUFDIR_wire\;
    \SIZ_wire\ <= SIZ;
    \TS_CPUn_wire\ <= TS_CPUn;
    CLKRAMA <= \CLKRAMA_wire\;
    TCI_CPUn <= \TCI_CPUn_wire\;
    CLKRAMB <= \CLKRAMB_wire\;
    BUFENn <= \BUFENn_wire\;
    \RnW_wire\ <= RnW;
    DMAn <= \DMAn_wire\;
    CLK80_CPU <= \CLK80_CPU_wire\;
    TSn <= \TSn_wire\;
    \PORTSIZE_wire\ <= PORTSIZE;
    \RESETn_wire\ <= RESETn;
    CLK40C <= \CLK40C_wire\;
    \BGn_wire\ <= BGn;
    TBI_CPUn <= \TBI_CPUn_wire\;
    CLK40A <= \CLK40A_wire\;
    \pll_pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll_pll\ : PLL40_2F
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            SCLK => '0',
            PLLOUTGLOBALA => \CLK80\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALB => \CLK40\,
            SDI => '0',
            PLLOUTCOREA => OPEN,
            BYPASS => '0',
            RESETB => \N__2891\,
            PLLOUTCOREB => OPEN,
            LOCK => OPEN,
            SDO => OPEN,
            EXTFEEDBACK => '0',
            DYNAMICDELAY => \pll_pll_DYNAMICDELAY_wire\,
            PLLIN => \N__8184\
        );

    \pll_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \VCCG0\,
            DIN => '0',
            DOUT => \N__8184\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \LBENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8168\,
            DIN => \N__8167\,
            DOUT => \N__8166\,
            PACKAGEPIN => \LBENn_wire\
        );

    \LBENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8168\,
            PADOUT => \N__8167\,
            PADIN => \N__8166\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \LBENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8159\,
            DIN => \N__8158\,
            DOUT => \N__8157\,
            PACKAGEPIN => D_UM_040(3)
        );

    \D_UM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8159\,
            PADOUT => \N__8158\,
            PADIN => \N__8157\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5417\,
            DIN0 => \D_UM_040_in_3\,
            DOUT0 => \N__7066\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TAn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8150\,
            DIN => \N__8149\,
            DOUT => \N__8148\,
            PACKAGEPIN => TAn
        );

    \TAn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8150\,
            PADOUT => \N__8149\,
            PADIN => \N__8148\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5788\,
            DIN0 => \TAn_in\,
            DOUT0 => \N__6316\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8141\,
            DIN => \N__8140\,
            DOUT => \N__8139\,
            PACKAGEPIN => D_LL_AMIGA(1)
        );

    \D_LL_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8141\,
            PADOUT => \N__8140\,
            PADIN => \N__8139\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2572\,
            DIN0 => \D_LL_AMIGA_in_1\,
            DOUT0 => \N__3898\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8132\,
            DIN => \N__8131\,
            DOUT => \N__8130\,
            PACKAGEPIN => D_UU_AMIGA(5)
        );

    \D_UU_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8132\,
            PADOUT => \N__8131\,
            PADIN => \N__8130\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2396\,
            DIN0 => \D_UU_AMIGA_in_5\,
            DOUT0 => \N__4084\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8123\,
            DIN => \N__8122\,
            DOUT => \N__8121\,
            PACKAGEPIN => D_UU_040(6)
        );

    \D_UU_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8123\,
            PADOUT => \N__8122\,
            PADIN => \N__8121\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5385\,
            DIN0 => \D_UU_040_in_6\,
            DOUT0 => \N__6520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUBGn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8114\,
            DIN => \N__8113\,
            DOUT => \N__8112\,
            PACKAGEPIN => \CPUBGn_wire\
        );

    \CPUBGn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8114\,
            PADOUT => \N__8113\,
            PADIN => \N__8112\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8105\,
            DIN => \N__8104\,
            DOUT => \N__8103\,
            PACKAGEPIN => D_LL_040(7)
        );

    \D_LL_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8105\,
            PADOUT => \N__8104\,
            PADIN => \N__8103\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5423\,
            DIN0 => \D_LL_040_in_7\,
            DOUT0 => \N__4336\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8096\,
            DIN => \N__8095\,
            DOUT => \N__8094\,
            PACKAGEPIN => D_LL_AMIGA(4)
        );

    \D_LL_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8096\,
            PADOUT => \N__8095\,
            PADIN => \N__8094\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2449\,
            DIN0 => \D_LL_AMIGA_in_4\,
            DOUT0 => \N__4215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8087\,
            DIN => \N__8086\,
            DOUT => \N__8085\,
            PACKAGEPIN => D_UM_AMIGA(3)
        );

    \D_UM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8087\,
            PADOUT => \N__8086\,
            PADIN => \N__8085\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2468\,
            DIN0 => \D_UM_AMIGA_in_3\,
            DOUT0 => \N__2917\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8078\,
            DIN => \N__8077\,
            DOUT => \N__8076\,
            PACKAGEPIN => D_UU_040(3)
        );

    \D_UU_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8078\,
            PADOUT => \N__8077\,
            PADIN => \N__8076\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5419\,
            DIN0 => \D_UU_040_in_3\,
            DOUT0 => \N__6655\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TEA_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8069\,
            DIN => \N__8068\,
            DOUT => \N__8067\,
            PACKAGEPIN => \TEA_CPUn_wire\
        );

    \TEA_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8069\,
            PADOUT => \N__8068\,
            PADIN => \N__8067\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2892\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8060\,
            DIN => \N__8059\,
            DOUT => \N__8058\,
            PACKAGEPIN => \A_040_wire\(1)
        );

    \A_040_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8060\,
            PADOUT => \N__8059\,
            PADIN => \N__8058\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8051\,
            DIN => \N__8050\,
            DOUT => \N__8049\,
            PACKAGEPIN => D_LM_AMIGA(3)
        );

    \D_LM_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8051\,
            PADOUT => \N__8050\,
            PADIN => \N__8049\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2531\,
            DIN0 => \D_LM_AMIGA_in_3\,
            DOUT0 => \N__4657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8042\,
            DIN => \N__8041\,
            DOUT => \N__8040\,
            PACKAGEPIN => D_LM_040(0)
        );

    \D_LM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8042\,
            PADOUT => \N__8041\,
            PADIN => \N__8040\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5424\,
            DIN0 => \D_LM_040_in_0\,
            DOUT0 => \N__4372\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8033\,
            DIN => \N__8032\,
            DOUT => \N__8031\,
            PACKAGEPIN => D_UM_AMIGA(6)
        );

    \D_UM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8033\,
            PADOUT => \N__8032\,
            PADIN => \N__8031\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2395\,
            DIN0 => \D_UM_AMIGA_in_6\,
            DOUT0 => \N__3142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8024\,
            DIN => \N__8023\,
            DOUT => \N__8022\,
            PACKAGEPIN => D_LM_AMIGA(4)
        );

    \D_LM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8024\,
            PADOUT => \N__8023\,
            PADIN => \N__8022\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2512\,
            DIN0 => \D_LM_AMIGA_in_4\,
            DOUT0 => \N__3727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8015\,
            DIN => \N__8014\,
            DOUT => \N__8013\,
            PACKAGEPIN => \A_AMIGA_wire\(1)
        );

    \A_AMIGA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8015\,
            PADOUT => \N__8014\,
            PADIN => \N__8013\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3915\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8006\,
            DIN => \N__8005\,
            DOUT => \N__8004\,
            PACKAGEPIN => D_LM_040(7)
        );

    \D_LM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__8006\,
            PADOUT => \N__8005\,
            PADIN => \N__8004\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5322\,
            DIN0 => \D_LM_040_in_7\,
            DOUT0 => \N__5002\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7997\,
            DIN => \N__7996\,
            DOUT => \N__7995\,
            PACKAGEPIN => D_UM_040(4)
        );

    \D_UM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7997\,
            PADOUT => \N__7996\,
            PADIN => \N__7995\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5420\,
            DIN0 => \D_UM_040_in_4\,
            DOUT0 => \N__7144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7988\,
            DIN => \N__7987\,
            DOUT => \N__7986\,
            PACKAGEPIN => \CLK40B_wire\
        );

    \CLK40B_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7988\,
            PADOUT => \N__7987\,
            PADIN => \N__7986\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4521\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7979\,
            DIN => \N__7978\,
            DOUT => \N__7977\,
            PACKAGEPIN => D_UU_AMIGA(0)
        );

    \D_UU_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7979\,
            PADOUT => \N__7978\,
            PADIN => \N__7977\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2475\,
            DIN0 => \D_UU_AMIGA_in_0\,
            DOUT0 => \N__2698\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7970\,
            DIN => \N__7969\,
            DOUT => \N__7968\,
            PACKAGEPIN => D_UM_040(1)
        );

    \D_UM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7970\,
            PADOUT => \N__7969\,
            PADIN => \N__7968\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5352\,
            DIN0 => \D_UM_040_in_1\,
            DOUT0 => \N__5719\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7961\,
            DIN => \N__7960\,
            DOUT => \N__7959\,
            PACKAGEPIN => D_LL_040(4)
        );

    \D_LL_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7961\,
            PADOUT => \N__7960\,
            PADIN => \N__7959\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5461\,
            DIN0 => \D_LL_040_in_4\,
            DOUT0 => \N__3538\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7952\,
            DIN => \N__7951\,
            DOUT => \N__7950\,
            PACKAGEPIN => D_LL_AMIGA(7)
        );

    \D_LL_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7952\,
            PADOUT => \N__7951\,
            PADIN => \N__7950\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2450\,
            DIN0 => \D_LL_AMIGA_in_7\,
            DOUT0 => \N__3430\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7943\,
            DIN => \N__7942\,
            DOUT => \N__7941\,
            PACKAGEPIN => D_UU_AMIGA(7)
        );

    \D_UU_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7943\,
            PADOUT => \N__7942\,
            PADIN => \N__7941\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2509\,
            DIN0 => \D_UU_AMIGA_in_7\,
            DOUT0 => \N__4003\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7934\,
            DIN => \N__7933\,
            DOUT => \N__7932\,
            PACKAGEPIN => \BUFDIR_wire\
        );

    \BUFDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7934\,
            PADOUT => \N__7933\,
            PADIN => \N__7932\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6052\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7925\,
            DIN => \N__7924\,
            DOUT => \N__7923\,
            PACKAGEPIN => D_LM_AMIGA(5)
        );

    \D_LM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7925\,
            PADOUT => \N__7924\,
            PADIN => \N__7923\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2488\,
            DIN0 => \D_LM_AMIGA_in_5\,
            DOUT0 => \N__4153\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7916\,
            DIN => \N__7915\,
            DOUT => \N__7914\,
            PACKAGEPIN => D_UU_040(4)
        );

    \D_UU_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7916\,
            PADOUT => \N__7915\,
            PADIN => \N__7914\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5381\,
            DIN0 => \D_UU_040_in_4\,
            DOUT0 => \N__6592\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7907\,
            DIN => \N__7906\,
            DOUT => \N__7905\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7907\,
            PADOUT => \N__7906\,
            PADIN => \N__7905\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7898\,
            DIN => \N__7897\,
            DOUT => \N__7896\,
            PACKAGEPIN => D_LM_040(6)
        );

    \D_LM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7898\,
            PADOUT => \N__7897\,
            PADIN => \N__7896\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5264\,
            DIN0 => \D_LM_040_in_6\,
            DOUT0 => \N__2995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7889\,
            DIN => \N__7888\,
            DOUT => \N__7887\,
            PACKAGEPIN => D_UM_040(5)
        );

    \D_UM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7889\,
            PADOUT => \N__7888\,
            PADIN => \N__7887\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5274\,
            DIN0 => \D_UM_040_in_5\,
            DOUT0 => \N__6718\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TS_CPUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7880\,
            DIN => \N__7879\,
            DOUT => \N__7878\,
            PACKAGEPIN => \TS_CPUn_wire\
        );

    \TS_CPUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7880\,
            PADOUT => \N__7879\,
            PADIN => \N__7878\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TS_CPUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7871\,
            DIN => \N__7870\,
            DOUT => \N__7869\,
            PACKAGEPIN => D_LL_040(1)
        );

    \D_LL_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7871\,
            PADOUT => \N__7870\,
            PADIN => \N__7869\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5452\,
            DIN0 => \D_LL_040_in_1\,
            DOUT0 => \N__3934\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7862\,
            DIN => \N__7861\,
            DOUT => \N__7860\,
            PACKAGEPIN => D_LL_AMIGA(3)
        );

    \D_LL_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7862\,
            PADOUT => \N__7861\,
            PADIN => \N__7860\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2573\,
            DIN0 => \D_LL_AMIGA_in_3\,
            DOUT0 => \N__2979\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7853\,
            DIN => \N__7852\,
            DOUT => \N__7851\,
            PACKAGEPIN => D_UM_AMIGA(5)
        );

    \D_UM_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7853\,
            PADOUT => \N__7852\,
            PADIN => \N__7851\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2508\,
            DIN0 => \D_UM_AMIGA_in_5\,
            DOUT0 => \N__4915\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7844\,
            DIN => \N__7843\,
            DOUT => \N__7842\,
            PACKAGEPIN => D_UU_040(1)
        );

    \D_UU_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7844\,
            PADOUT => \N__7843\,
            PADIN => \N__7842\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5418\,
            DIN0 => \D_UU_040_in_1\,
            DOUT0 => \N__5932\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7835\,
            DIN => \N__7834\,
            DOUT => \N__7833\,
            PACKAGEPIN => D_UU_AMIGA(3)
        );

    \D_UU_AMIGA_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7835\,
            PADOUT => \N__7834\,
            PADIN => \N__7833\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2511\,
            DIN0 => \D_UU_AMIGA_in_3\,
            DOUT0 => \N__4609\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7826\,
            DIN => \N__7825\,
            DOUT => \N__7824\,
            PACKAGEPIN => D_LM_AMIGA(1)
        );

    \D_LM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7826\,
            PADOUT => \N__7825\,
            PADIN => \N__7824\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2542\,
            DIN0 => \D_LM_AMIGA_in_1\,
            DOUT0 => \N__3799\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7817\,
            DIN => \N__7816\,
            DOUT => \N__7815\,
            PACKAGEPIN => D_LM_040(2)
        );

    \D_LM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7817\,
            PADOUT => \N__7816\,
            PADIN => \N__7815\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5422\,
            DIN0 => \D_LM_040_in_2\,
            DOUT0 => \N__3445\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7808\,
            DIN => \N__7807\,
            DOUT => \N__7806\,
            PACKAGEPIN => D_LL_040(5)
        );

    \D_LL_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7808\,
            PADOUT => \N__7807\,
            PADIN => \N__7806\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5425\,
            DIN0 => \D_LL_040_in_5\,
            DOUT0 => \N__3262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7799\,
            DIN => \N__7798\,
            DOUT => \N__7797\,
            PACKAGEPIN => D_LL_AMIGA(6)
        );

    \D_LL_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7799\,
            PADOUT => \N__7798\,
            PADIN => \N__7797\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2558\,
            DIN0 => \D_LL_AMIGA_in_6\,
            DOUT0 => \N__3187\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7790\,
            DIN => \N__7789\,
            DOUT => \N__7788\,
            PACKAGEPIN => D_UU_AMIGA(6)
        );

    \D_UU_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7790\,
            PADOUT => \N__7789\,
            PADIN => \N__7788\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2510\,
            DIN0 => \D_UU_AMIGA_in_6\,
            DOUT0 => \N__2785\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7781\,
            DIN => \N__7780\,
            DOUT => \N__7779\,
            PACKAGEPIN => D_UM_AMIGA(1)
        );

    \D_UM_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7781\,
            PADOUT => \N__7780\,
            PADIN => \N__7779\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2489\,
            DIN0 => \D_UM_AMIGA_in_1\,
            DOUT0 => \N__3838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7772\,
            DIN => \N__7771\,
            DOUT => \N__7770\,
            PACKAGEPIN => D_UU_040(5)
        );

    \D_UU_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7772\,
            PADOUT => \N__7771\,
            PADIN => \N__7770\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5275\,
            DIN0 => \D_UU_040_in_5\,
            DOUT0 => \N__6799\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7763\,
            DIN => \N__7762\,
            DOUT => \N__7761\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7763\,
            PADOUT => \N__7762\,
            PADIN => \N__7761\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__3301\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__2644\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7754\,
            DIN => \N__7753\,
            DOUT => \N__7752\,
            PACKAGEPIN => \CLKRAMA_wire\
        );

    \CLKRAMA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7754\,
            PADOUT => \N__7753\,
            PADIN => \N__7752\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4525\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7745\,
            DIN => \N__7744\,
            DOUT => \N__7743\,
            PACKAGEPIN => D_UM_040(2)
        );

    \D_UM_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7745\,
            PADOUT => \N__7744\,
            PADIN => \N__7743\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5313\,
            DIN0 => \D_UM_040_in_2\,
            DOUT0 => \N__6499\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7736\,
            DIN => \N__7735\,
            DOUT => \N__7734\,
            PACKAGEPIN => D_LL_040(2)
        );

    \D_LL_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7736\,
            PADOUT => \N__7735\,
            PADIN => \N__7734\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5439\,
            DIN0 => \D_LL_040_in_2\,
            DOUT0 => \N__3568\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7727\,
            DIN => \N__7726\,
            DOUT => \N__7725\,
            PACKAGEPIN => \TCI_CPUn_wire\
        );

    \TCI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7727\,
            PADOUT => \N__7726\,
            PADIN => \N__7725\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2882\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAMB_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7718\,
            DIN => \N__7717\,
            DOUT => \N__7716\,
            PACKAGEPIN => \CLKRAMB_wire\
        );

    \CLKRAMB_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7718\,
            PADOUT => \N__7717\,
            PADIN => \N__7716\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7709\,
            DIN => \N__7708\,
            DOUT => \N__7707\,
            PACKAGEPIN => D_LL_AMIGA(2)
        );

    \D_LL_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7709\,
            PADOUT => \N__7708\,
            PADIN => \N__7707\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2574\,
            DIN0 => \D_LL_AMIGA_in_2\,
            DOUT0 => \N__3121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7700\,
            DIN => \N__7699\,
            DOUT => \N__7698\,
            PACKAGEPIN => D_UM_AMIGA(4)
        );

    \D_UM_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7700\,
            PADOUT => \N__7699\,
            PADIN => \N__7698\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2472\,
            DIN0 => \D_UM_AMIGA_in_4\,
            DOUT0 => \N__4168\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7691\,
            DIN => \N__7690\,
            DOUT => \N__7689\,
            PACKAGEPIN => D_UU_AMIGA(2)
        );

    \D_UU_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7691\,
            PADOUT => \N__7690\,
            PADIN => \N__7689\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2474\,
            DIN0 => \D_UU_AMIGA_in_2\,
            DOUT0 => \N__3604\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7682\,
            DIN => \N__7681\,
            DOUT => \N__7680\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7682\,
            PADOUT => \N__7681\,
            PADIN => \N__7680\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3820\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7673\,
            DIN => \N__7672\,
            DOUT => \N__7671\,
            PACKAGEPIN => D_LM_AMIGA(6)
        );

    \D_LM_AMIGA_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7673\,
            PADOUT => \N__7672\,
            PADIN => \N__7671\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2453\,
            DIN0 => \D_LM_AMIGA_in_6\,
            DOUT0 => \N__2821\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7664\,
            DIN => \N__7663\,
            DOUT => \N__7662\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7664\,
            PADOUT => \N__7663\,
            PADIN => \N__7662\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7655\,
            DIN => \N__7654\,
            DOUT => \N__7653\,
            PACKAGEPIN => D_LM_040(5)
        );

    \D_LM_040_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7655\,
            PADOUT => \N__7654\,
            PADIN => \N__7653\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5331\,
            DIN0 => \D_LM_040_in_5\,
            DOUT0 => \N__3037\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7646\,
            DIN => \N__7645\,
            DOUT => \N__7644\,
            PACKAGEPIN => D_UM_040(6)
        );

    \D_UM_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7646\,
            PADOUT => \N__7645\,
            PADIN => \N__7644\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5224\,
            DIN0 => \D_UM_040_in_6\,
            DOUT0 => \N__6481\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMAn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7637\,
            DIN => \N__7636\,
            DOUT => \N__7635\,
            PACKAGEPIN => \DMAn_wire\
        );

    \DMAn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7637\,
            PADOUT => \N__7636\,
            PADIN => \N__7635\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2896\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7628\,
            DIN => \N__7627\,
            DOUT => \N__7626\,
            PACKAGEPIN => D_LL_040(6)
        );

    \D_LL_040_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7628\,
            PADOUT => \N__7627\,
            PADIN => \N__7626\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5426\,
            DIN0 => \D_LL_040_in_6\,
            DOUT0 => \N__3502\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7619\,
            DIN => \N__7618\,
            DOUT => \N__7617\,
            PACKAGEPIN => D_LL_AMIGA(5)
        );

    \D_LL_AMIGA_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7619\,
            PADOUT => \N__7618\,
            PADIN => \N__7617\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2559\,
            DIN0 => \D_LL_AMIGA_in_5\,
            DOUT0 => \N__4984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7610\,
            DIN => \N__7609\,
            DOUT => \N__7608\,
            PACKAGEPIN => D_UM_AMIGA(0)
        );

    \D_UM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7610\,
            PADOUT => \N__7609\,
            PADIN => \N__7608\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2530\,
            DIN0 => \D_UM_AMIGA_in_0\,
            DOUT0 => \N__4258\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7601\,
            DIN => \N__7600\,
            DOUT => \N__7599\,
            PACKAGEPIN => D_UU_040(2)
        );

    \D_UU_040_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7601\,
            PADOUT => \N__7600\,
            PADIN => \N__7599\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5382\,
            DIN0 => \D_UU_040_in_2\,
            DOUT0 => \N__5512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7592\,
            DIN => \N__7591\,
            DOUT => \N__7590\,
            PACKAGEPIN => D_LM_AMIGA(2)
        );

    \D_LM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7592\,
            PADOUT => \N__7591\,
            PADIN => \N__7590\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2529\,
            DIN0 => \D_LM_AMIGA_in_2\,
            DOUT0 => \N__3636\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK80_CPU_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7583\,
            DIN => \N__7582\,
            DOUT => \N__7581\,
            PACKAGEPIN => \CLK80_CPU_wire\
        );

    \CLK80_CPU_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7583\,
            PADOUT => \N__7582\,
            PADIN => \N__7581\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4422\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7574\,
            DIN => \N__7573\,
            DOUT => \N__7572\,
            PACKAGEPIN => D_LL_040(3)
        );

    \D_LL_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7574\,
            PADOUT => \N__7573\,
            PADIN => \N__7572\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5456\,
            DIN0 => \D_LL_040_in_3\,
            DOUT0 => \N__3970\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7565\,
            DIN => \N__7564\,
            DOUT => \N__7563\,
            PACKAGEPIN => D_LM_040(1)
        );

    \D_LM_040_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7565\,
            PADOUT => \N__7564\,
            PADIN => \N__7563\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5421\,
            DIN0 => \D_LM_040_in_1\,
            DOUT0 => \N__4543\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7556\,
            DIN => \N__7555\,
            DOUT => \N__7554\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7556\,
            PADOUT => \N__7555\,
            PADIN => \N__7554\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3292\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7547\,
            DIN => \N__7546\,
            DOUT => \N__7545\,
            PACKAGEPIN => D_UM_AMIGA(7)
        );

    \D_UM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7547\,
            PADOUT => \N__7546\,
            PADIN => \N__7545\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2507\,
            DIN0 => \D_UM_AMIGA_in_7\,
            DOUT0 => \N__3364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7538\,
            DIN => \N__7537\,
            DOUT => \N__7536\,
            PACKAGEPIN => D_LM_AMIGA(7)
        );

    \D_LM_AMIGA_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7538\,
            PADOUT => \N__7537\,
            PADIN => \N__7536\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2452\,
            DIN0 => \D_LM_AMIGA_in_7\,
            DOUT0 => \N__4063\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7529\,
            DIN => \N__7528\,
            DOUT => \N__7527\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7529\,
            PADOUT => \N__7528\,
            PADIN => \N__7527\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PORTSIZE_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_AMIGA_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7520\,
            DIN => \N__7519\,
            DOUT => \N__7518\,
            PACKAGEPIN => \A_AMIGA_wire\(0)
        );

    \A_AMIGA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7520\,
            PADOUT => \N__7519\,
            PADIN => \N__7518\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7511\,
            DIN => \N__7510\,
            DOUT => \N__7509\,
            PACKAGEPIN => D_LM_040(4)
        );

    \D_LM_040_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7511\,
            PADOUT => \N__7510\,
            PADIN => \N__7509\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5353\,
            DIN0 => \D_LM_040_in_4\,
            DOUT0 => \N__3223\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7502\,
            DIN => \N__7501\,
            DOUT => \N__7500\,
            PACKAGEPIN => D_UM_040(7)
        );

    \D_UM_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7502\,
            PADOUT => \N__7501\,
            PADIN => \N__7500\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5416\,
            DIN0 => \D_UM_040_in_7\,
            DOUT0 => \N__6931\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7493\,
            DIN => \N__7492\,
            DOUT => \N__7491\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7493\,
            PADOUT => \N__7492\,
            PADIN => \N__7491\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7484\,
            DIN => \N__7483\,
            DOUT => \N__7482\,
            PACKAGEPIN => D_UU_AMIGA(1)
        );

    \D_UU_AMIGA_iobuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7484\,
            PADOUT => \N__7483\,
            PADIN => \N__7482\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2467\,
            DIN0 => \D_UU_AMIGA_in_1\,
            DOUT0 => \N__3742\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7475\,
            DIN => \N__7474\,
            DOUT => \N__7473\,
            PACKAGEPIN => \CLK40C_wire\
        );

    \CLK40C_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7475\,
            PADOUT => \N__7474\,
            PADIN => \N__7473\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7466\,
            DIN => \N__7465\,
            DOUT => \N__7464\,
            PACKAGEPIN => D_UM_040(0)
        );

    \D_UM_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7466\,
            PADOUT => \N__7465\,
            PADIN => \N__7464\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5330\,
            DIN0 => \D_UM_040_in_0\,
            DOUT0 => \N__5500\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7457\,
            DIN => \N__7456\,
            DOUT => \N__7455\,
            PACKAGEPIN => D_LL_AMIGA(0)
        );

    \D_LL_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7457\,
            PADOUT => \N__7456\,
            PADIN => \N__7455\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2578\,
            DIN0 => \D_LL_AMIGA_in_0\,
            DOUT0 => \N__4315\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_AMIGA_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7448\,
            DIN => \N__7447\,
            DOUT => \N__7446\,
            PACKAGEPIN => D_UU_AMIGA(4)
        );

    \D_UU_AMIGA_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7448\,
            PADOUT => \N__7447\,
            PADIN => \N__7446\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2473\,
            DIN0 => \D_UU_AMIGA_in_4\,
            DOUT0 => \N__3673\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7439\,
            DIN => \N__7438\,
            DOUT => \N__7437\,
            PACKAGEPIN => D_UU_040(7)
        );

    \D_UU_040_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7439\,
            PADOUT => \N__7438\,
            PADIN => \N__7437\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5384\,
            DIN0 => \D_UU_040_in_7\,
            DOUT0 => \N__5578\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7430\,
            DIN => \N__7429\,
            DOUT => \N__7428\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7430\,
            PADOUT => \N__7429\,
            PADIN => \N__7428\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BGn_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7421\,
            DIN => \N__7420\,
            DOUT => \N__7419\,
            PACKAGEPIN => \BGn_wire\
        );

    \BGn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7421\,
            PADOUT => \N__7420\,
            PADIN => \N__7419\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \BGn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LL_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7412\,
            DIN => \N__7411\,
            DOUT => \N__7410\,
            PACKAGEPIN => D_LL_040(0)
        );

    \D_LL_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7412\,
            PADOUT => \N__7411\,
            PADIN => \N__7410\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5457\,
            DIN0 => \D_LL_040_in_0\,
            DOUT0 => \N__3325\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UM_AMIGA_iobuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7403\,
            DIN => \N__7402\,
            DOUT => \N__7401\,
            PACKAGEPIN => D_UM_AMIGA(2)
        );

    \D_UM_AMIGA_iobuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7403\,
            PADOUT => \N__7402\,
            PADIN => \N__7401\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2513\,
            DIN0 => \D_UM_AMIGA_in_2\,
            DOUT0 => \N__3070\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_UU_040_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7394\,
            DIN => \N__7393\,
            DOUT => \N__7392\,
            PACKAGEPIN => D_UU_040(0)
        );

    \D_UU_040_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7394\,
            PADOUT => \N__7393\,
            PADIN => \N__7392\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5383\,
            DIN0 => \D_UU_040_in_0\,
            DOUT0 => \N__6868\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_040_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__7385\,
            DIN => \N__7384\,
            DOUT => \N__7383\,
            PACKAGEPIN => \A_040_wire\(0)
        );

    \A_040_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7385\,
            PADOUT => \N__7384\,
            PADIN => \N__7383\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_040_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_AMIGA_iobuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7376\,
            DIN => \N__7375\,
            DOUT => \N__7374\,
            PACKAGEPIN => D_LM_AMIGA(0)
        );

    \D_LM_AMIGA_iobuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7376\,
            PADOUT => \N__7375\,
            PADIN => \N__7374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__2451\,
            DIN0 => \D_LM_AMIGA_in_0\,
            DOUT0 => \N__2746\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBI_CPUn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7367\,
            DIN => \N__7366\,
            DOUT => \N__7365\,
            PACKAGEPIN => \TBI_CPUn_wire\
        );

    \TBI_CPUn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7367\,
            PADOUT => \N__7366\,
            PADIN => \N__7365\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4585\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40A_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7358\,
            DIN => \N__7357\,
            DOUT => \N__7356\,
            PACKAGEPIN => \CLK40A_wire\
        );

    \CLK40A_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7358\,
            PADOUT => \N__7357\,
            PADIN => \N__7356\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4519\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_LM_040_iobuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7349\,
            DIN => \N__7348\,
            DOUT => \N__7347\,
            PACKAGEPIN => D_LM_040(3)
        );

    \D_LM_040_iobuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__7349\,
            PADOUT => \N__7348\,
            PADIN => \N__7347\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5392\,
            DIN0 => \D_LM_040_in_3\,
            DOUT0 => \N__2665\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1874\ : InMux
    port map (
            O => \N__7330\,
            I => \N__7327\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\
        );

    \I__1872\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7321\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__7321\,
            I => \N__7316\
        );

    \I__1870\ : InMux
    port map (
            O => \N__7320\,
            I => \N__7313\
        );

    \I__1869\ : InMux
    port map (
            O => \N__7319\,
            I => \N__7310\
        );

    \I__1868\ : Span4Mux_v
    port map (
            O => \N__7316\,
            I => \N__7307\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__7313\,
            I => \N__7302\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__7310\,
            I => \N__7302\
        );

    \I__1865\ : Span4Mux_v
    port map (
            O => \N__7307\,
            I => \N__7299\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__7302\,
            I => \N__7296\
        );

    \I__1863\ : Sp12to4
    port map (
            O => \N__7299\,
            I => \N__7293\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__7296\,
            I => \N__7290\
        );

    \I__1861\ : Span12Mux_h
    port map (
            O => \N__7293\,
            I => \N__7287\
        );

    \I__1860\ : Sp12to4
    port map (
            O => \N__7290\,
            I => \N__7284\
        );

    \I__1859\ : Span12Mux_v
    port map (
            O => \N__7287\,
            I => \N__7281\
        );

    \I__1858\ : Span12Mux_h
    port map (
            O => \N__7284\,
            I => \N__7278\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__7281\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1856\ : Odrv12
    port map (
            O => \N__7278\,
            I => \D_UM_AMIGA_in_4\
        );

    \I__1855\ : InMux
    port map (
            O => \N__7273\,
            I => \N__7267\
        );

    \I__1854\ : InMux
    port map (
            O => \N__7272\,
            I => \N__7267\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__7267\,
            I => \N__7264\
        );

    \I__1852\ : Span4Mux_v
    port map (
            O => \N__7264\,
            I => \N__7254\
        );

    \I__1851\ : InMux
    port map (
            O => \N__7263\,
            I => \N__7251\
        );

    \I__1850\ : InMux
    port map (
            O => \N__7262\,
            I => \N__7243\
        );

    \I__1849\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7243\
        );

    \I__1848\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7234\
        );

    \I__1847\ : InMux
    port map (
            O => \N__7259\,
            I => \N__7234\
        );

    \I__1846\ : InMux
    port map (
            O => \N__7258\,
            I => \N__7234\
        );

    \I__1845\ : InMux
    port map (
            O => \N__7257\,
            I => \N__7234\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__7254\,
            I => \N__7224\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__7251\,
            I => \N__7221\
        );

    \I__1842\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7216\
        );

    \I__1841\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7216\
        );

    \I__1840\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7213\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__7243\,
            I => \N__7210\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__7234\,
            I => \N__7207\
        );

    \I__1837\ : InMux
    port map (
            O => \N__7233\,
            I => \N__7200\
        );

    \I__1836\ : InMux
    port map (
            O => \N__7232\,
            I => \N__7200\
        );

    \I__1835\ : InMux
    port map (
            O => \N__7231\,
            I => \N__7200\
        );

    \I__1834\ : InMux
    port map (
            O => \N__7230\,
            I => \N__7195\
        );

    \I__1833\ : InMux
    port map (
            O => \N__7229\,
            I => \N__7195\
        );

    \I__1832\ : InMux
    port map (
            O => \N__7228\,
            I => \N__7190\
        );

    \I__1831\ : InMux
    port map (
            O => \N__7227\,
            I => \N__7190\
        );

    \I__1830\ : Span12Mux_h
    port map (
            O => \N__7224\,
            I => \N__7185\
        );

    \I__1829\ : Span4Mux_h
    port map (
            O => \N__7221\,
            I => \N__7180\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__7216\,
            I => \N__7180\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__7213\,
            I => \N__7177\
        );

    \I__1826\ : Span4Mux_v
    port map (
            O => \N__7210\,
            I => \N__7170\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__7207\,
            I => \N__7170\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__7200\,
            I => \N__7170\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__7195\,
            I => \N__7165\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__7190\,
            I => \N__7165\
        );

    \I__1821\ : InMux
    port map (
            O => \N__7189\,
            I => \N__7162\
        );

    \I__1820\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7159\
        );

    \I__1819\ : Odrv12
    port map (
            O => \N__7185\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__7180\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__7177\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__7170\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1815\ : Odrv12
    port map (
            O => \N__7165\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__7162\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__7159\,
            I => \U111_CYCLE_SM.LW_CYCLEZ0\
        );

    \I__1812\ : IoInMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1810\ : IoSpan4Mux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1809\ : Span4Mux_s3_v
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1808\ : Sp12to4
    port map (
            O => \N__7132\,
            I => \N__7129\
        );

    \I__1807\ : Span12Mux_h
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1806\ : Odrv12
    port map (
            O => \N__7126\,
            I => \un1_D_UM_AMIGA_4\
        );

    \I__1805\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7120\
        );

    \I__1804\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7116\
        );

    \I__1803\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7113\
        );

    \I__1802\ : Span4Mux_v
    port map (
            O => \N__7116\,
            I => \N__7109\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__7113\,
            I => \N__7106\
        );

    \I__1800\ : InMux
    port map (
            O => \N__7112\,
            I => \N__7103\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__7109\,
            I => \N__7100\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__7106\,
            I => \N__7095\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7103\,
            I => \N__7095\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__7100\,
            I => \N__7092\
        );

    \I__1795\ : Span4Mux_v
    port map (
            O => \N__7095\,
            I => \N__7089\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__7092\,
            I => \N__7086\
        );

    \I__1793\ : Sp12to4
    port map (
            O => \N__7089\,
            I => \N__7083\
        );

    \I__1792\ : Span12Mux_v
    port map (
            O => \N__7086\,
            I => \N__7078\
        );

    \I__1791\ : Span12Mux_h
    port map (
            O => \N__7083\,
            I => \N__7078\
        );

    \I__1790\ : Odrv12
    port map (
            O => \N__7078\,
            I => \D_UM_AMIGA_in_3\
        );

    \I__1789\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7072\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1787\ : Odrv12
    port map (
            O => \N__7069\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\
        );

    \I__1786\ : IoInMux
    port map (
            O => \N__7066\,
            I => \N__7063\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__7063\,
            I => \N__7060\
        );

    \I__1784\ : IoSpan4Mux
    port map (
            O => \N__7060\,
            I => \N__7057\
        );

    \I__1783\ : IoSpan4Mux
    port map (
            O => \N__7057\,
            I => \N__7054\
        );

    \I__1782\ : Span4Mux_s2_h
    port map (
            O => \N__7054\,
            I => \N__7051\
        );

    \I__1781\ : Sp12to4
    port map (
            O => \N__7051\,
            I => \N__7048\
        );

    \I__1780\ : Odrv12
    port map (
            O => \N__7048\,
            I => \un1_D_UM_AMIGA_3\
        );

    \I__1779\ : CEMux
    port map (
            O => \N__7045\,
            I => \N__7040\
        );

    \I__1778\ : CEMux
    port map (
            O => \N__7044\,
            I => \N__7037\
        );

    \I__1777\ : CEMux
    port map (
            O => \N__7043\,
            I => \N__7033\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__7040\,
            I => \N__7028\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__7037\,
            I => \N__7028\
        );

    \I__1774\ : CEMux
    port map (
            O => \N__7036\,
            I => \N__7025\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__7033\,
            I => \N__7022\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__7028\,
            I => \N__7017\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__7025\,
            I => \N__7017\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__7022\,
            I => \N__7014\
        );

    \I__1769\ : Span4Mux_h
    port map (
            O => \N__7017\,
            I => \N__7011\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__7014\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1767\ : Odrv4
    port map (
            O => \N__7011\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\
        );

    \I__1766\ : SRMux
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__1765\ : SRMux
    port map (
            O => \N__7005\,
            I => \N__6997\
        );

    \I__1764\ : SRMux
    port map (
            O => \N__7004\,
            I => \N__6994\
        );

    \I__1763\ : SRMux
    port map (
            O => \N__7003\,
            I => \N__6991\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7000\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__6997\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__6994\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__6991\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\
        );

    \I__1758\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6979\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__6979\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\
        );

    \I__1756\ : InMux
    port map (
            O => \N__6976\,
            I => \N__6971\
        );

    \I__1755\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6968\
        );

    \I__1754\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6965\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__6971\,
            I => \N__6960\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__6968\,
            I => \N__6960\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__6965\,
            I => \N__6957\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__6960\,
            I => \N__6954\
        );

    \I__1749\ : Span12Mux_v
    port map (
            O => \N__6957\,
            I => \N__6951\
        );

    \I__1748\ : Span4Mux_v
    port map (
            O => \N__6954\,
            I => \N__6948\
        );

    \I__1747\ : Span12Mux_h
    port map (
            O => \N__6951\,
            I => \N__6945\
        );

    \I__1746\ : Sp12to4
    port map (
            O => \N__6948\,
            I => \N__6942\
        );

    \I__1745\ : Span12Mux_v
    port map (
            O => \N__6945\,
            I => \N__6939\
        );

    \I__1744\ : Span12Mux_h
    port map (
            O => \N__6942\,
            I => \N__6936\
        );

    \I__1743\ : Odrv12
    port map (
            O => \N__6939\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1742\ : Odrv12
    port map (
            O => \N__6936\,
            I => \D_UM_AMIGA_in_7\
        );

    \I__1741\ : IoInMux
    port map (
            O => \N__6931\,
            I => \N__6928\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__6928\,
            I => \N__6925\
        );

    \I__1739\ : Sp12to4
    port map (
            O => \N__6925\,
            I => \N__6922\
        );

    \I__1738\ : Span12Mux_h
    port map (
            O => \N__6922\,
            I => \N__6919\
        );

    \I__1737\ : Odrv12
    port map (
            O => \N__6919\,
            I => \un1_D_UM_AMIGA_7\
        );

    \I__1736\ : InMux
    port map (
            O => \N__6916\,
            I => \N__6913\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__6913\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\
        );

    \I__1734\ : InMux
    port map (
            O => \N__6910\,
            I => \N__6907\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__6907\,
            I => \N__6902\
        );

    \I__1732\ : InMux
    port map (
            O => \N__6906\,
            I => \N__6899\
        );

    \I__1731\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6896\
        );

    \I__1730\ : Span4Mux_v
    port map (
            O => \N__6902\,
            I => \N__6893\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__6899\,
            I => \N__6888\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__6896\,
            I => \N__6888\
        );

    \I__1727\ : Span4Mux_v
    port map (
            O => \N__6893\,
            I => \N__6885\
        );

    \I__1726\ : Span4Mux_v
    port map (
            O => \N__6888\,
            I => \N__6882\
        );

    \I__1725\ : Span4Mux_v
    port map (
            O => \N__6885\,
            I => \N__6877\
        );

    \I__1724\ : Span4Mux_h
    port map (
            O => \N__6882\,
            I => \N__6877\
        );

    \I__1723\ : Sp12to4
    port map (
            O => \N__6877\,
            I => \N__6874\
        );

    \I__1722\ : Span12Mux_h
    port map (
            O => \N__6874\,
            I => \N__6871\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__6871\,
            I => \D_UU_AMIGA_in_0\
        );

    \I__1720\ : IoInMux
    port map (
            O => \N__6868\,
            I => \N__6865\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6862\
        );

    \I__1718\ : Span4Mux_s3_v
    port map (
            O => \N__6862\,
            I => \N__6859\
        );

    \I__1717\ : Span4Mux_h
    port map (
            O => \N__6859\,
            I => \N__6856\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__6856\,
            I => \N__6853\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__6853\,
            I => \N__6850\
        );

    \I__1714\ : Odrv4
    port map (
            O => \N__6850\,
            I => \un1_D_UU_AMIGA_0\
        );

    \I__1713\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__6844\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\
        );

    \I__1711\ : InMux
    port map (
            O => \N__6841\,
            I => \N__6838\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__6838\,
            I => \N__6834\
        );

    \I__1709\ : InMux
    port map (
            O => \N__6837\,
            I => \N__6831\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__6834\,
            I => \N__6826\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__6831\,
            I => \N__6826\
        );

    \I__1706\ : Span4Mux_h
    port map (
            O => \N__6826\,
            I => \N__6822\
        );

    \I__1705\ : InMux
    port map (
            O => \N__6825\,
            I => \N__6819\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__6822\,
            I => \N__6814\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__6819\,
            I => \N__6814\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1701\ : Sp12to4
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__1700\ : Span12Mux_h
    port map (
            O => \N__6808\,
            I => \N__6805\
        );

    \I__1699\ : Span12Mux_v
    port map (
            O => \N__6805\,
            I => \N__6802\
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__6802\,
            I => \D_UU_AMIGA_in_5\
        );

    \I__1697\ : IoInMux
    port map (
            O => \N__6799\,
            I => \N__6796\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__6796\,
            I => \N__6793\
        );

    \I__1695\ : Span4Mux_s3_v
    port map (
            O => \N__6793\,
            I => \N__6790\
        );

    \I__1694\ : Span4Mux_v
    port map (
            O => \N__6790\,
            I => \N__6787\
        );

    \I__1693\ : Sp12to4
    port map (
            O => \N__6787\,
            I => \N__6784\
        );

    \I__1692\ : Span12Mux_h
    port map (
            O => \N__6784\,
            I => \N__6781\
        );

    \I__1691\ : Odrv12
    port map (
            O => \N__6781\,
            I => \un1_D_UU_AMIGA_5\
        );

    \I__1690\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6775\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__6775\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\
        );

    \I__1688\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6768\
        );

    \I__1687\ : InMux
    port map (
            O => \N__6771\,
            I => \N__6765\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__6768\,
            I => \N__6761\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__6765\,
            I => \N__6758\
        );

    \I__1684\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6755\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__6761\,
            I => \N__6752\
        );

    \I__1682\ : Span4Mux_v
    port map (
            O => \N__6758\,
            I => \N__6749\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6746\
        );

    \I__1680\ : Sp12to4
    port map (
            O => \N__6752\,
            I => \N__6743\
        );

    \I__1679\ : Sp12to4
    port map (
            O => \N__6749\,
            I => \N__6740\
        );

    \I__1678\ : Span12Mux_h
    port map (
            O => \N__6746\,
            I => \N__6737\
        );

    \I__1677\ : Span12Mux_h
    port map (
            O => \N__6743\,
            I => \N__6734\
        );

    \I__1676\ : Span12Mux_h
    port map (
            O => \N__6740\,
            I => \N__6731\
        );

    \I__1675\ : Span12Mux_h
    port map (
            O => \N__6737\,
            I => \N__6728\
        );

    \I__1674\ : Span12Mux_v
    port map (
            O => \N__6734\,
            I => \N__6723\
        );

    \I__1673\ : Span12Mux_h
    port map (
            O => \N__6731\,
            I => \N__6723\
        );

    \I__1672\ : Odrv12
    port map (
            O => \N__6728\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1671\ : Odrv12
    port map (
            O => \N__6723\,
            I => \D_UM_AMIGA_in_5\
        );

    \I__1670\ : IoInMux
    port map (
            O => \N__6718\,
            I => \N__6715\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__6715\,
            I => \N__6712\
        );

    \I__1668\ : Span4Mux_s2_v
    port map (
            O => \N__6712\,
            I => \N__6709\
        );

    \I__1667\ : Sp12to4
    port map (
            O => \N__6709\,
            I => \N__6706\
        );

    \I__1666\ : Span12Mux_h
    port map (
            O => \N__6706\,
            I => \N__6703\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__6703\,
            I => \un1_D_UM_AMIGA_5\
        );

    \I__1664\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6697\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__6697\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\
        );

    \I__1662\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6690\
        );

    \I__1661\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6687\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__6690\,
            I => \N__6684\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__6687\,
            I => \N__6681\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__6684\,
            I => \N__6675\
        );

    \I__1657\ : Span4Mux_v
    port map (
            O => \N__6681\,
            I => \N__6675\
        );

    \I__1656\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6672\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__6675\,
            I => \N__6667\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__6672\,
            I => \N__6667\
        );

    \I__1653\ : Sp12to4
    port map (
            O => \N__6667\,
            I => \N__6664\
        );

    \I__1652\ : Span12Mux_v
    port map (
            O => \N__6664\,
            I => \N__6661\
        );

    \I__1651\ : Span12Mux_h
    port map (
            O => \N__6661\,
            I => \N__6658\
        );

    \I__1650\ : Odrv12
    port map (
            O => \N__6658\,
            I => \D_UU_AMIGA_in_3\
        );

    \I__1649\ : IoInMux
    port map (
            O => \N__6655\,
            I => \N__6652\
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1647\ : Span12Mux_s0_v
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1646\ : Span12Mux_h
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__6643\,
            I => \un1_D_UU_AMIGA_3\
        );

    \I__1644\ : InMux
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__6637\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\
        );

    \I__1642\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6631\,
            I => \N__6626\
        );

    \I__1640\ : InMux
    port map (
            O => \N__6630\,
            I => \N__6623\
        );

    \I__1639\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6620\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__6626\,
            I => \N__6617\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__6623\,
            I => \N__6612\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__6620\,
            I => \N__6612\
        );

    \I__1635\ : Sp12to4
    port map (
            O => \N__6617\,
            I => \N__6609\
        );

    \I__1634\ : Span12Mux_v
    port map (
            O => \N__6612\,
            I => \N__6606\
        );

    \I__1633\ : Span12Mux_h
    port map (
            O => \N__6609\,
            I => \N__6603\
        );

    \I__1632\ : Span12Mux_h
    port map (
            O => \N__6606\,
            I => \N__6600\
        );

    \I__1631\ : Span12Mux_v
    port map (
            O => \N__6603\,
            I => \N__6597\
        );

    \I__1630\ : Odrv12
    port map (
            O => \N__6600\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1629\ : Odrv12
    port map (
            O => \N__6597\,
            I => \D_UU_AMIGA_in_4\
        );

    \I__1628\ : IoInMux
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1626\ : Span4Mux_s2_v
    port map (
            O => \N__6586\,
            I => \N__6583\
        );

    \I__1625\ : Span4Mux_h
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1623\ : Span4Mux_v
    port map (
            O => \N__6577\,
            I => \N__6574\
        );

    \I__1622\ : Odrv4
    port map (
            O => \N__6574\,
            I => \un1_D_UU_AMIGA_4\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__6568\,
            I => \N__6565\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__6565\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\
        );

    \I__1618\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6558\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6555\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__6558\,
            I => \N__6551\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__6555\,
            I => \N__6548\
        );

    \I__1614\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6545\
        );

    \I__1613\ : Span4Mux_v
    port map (
            O => \N__6551\,
            I => \N__6540\
        );

    \I__1612\ : Span4Mux_v
    port map (
            O => \N__6548\,
            I => \N__6540\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__6545\,
            I => \N__6537\
        );

    \I__1610\ : Span4Mux_h
    port map (
            O => \N__6540\,
            I => \N__6534\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__6537\,
            I => \N__6531\
        );

    \I__1608\ : Sp12to4
    port map (
            O => \N__6534\,
            I => \N__6526\
        );

    \I__1607\ : Sp12to4
    port map (
            O => \N__6531\,
            I => \N__6526\
        );

    \I__1606\ : Span12Mux_h
    port map (
            O => \N__6526\,
            I => \N__6523\
        );

    \I__1605\ : Odrv12
    port map (
            O => \N__6523\,
            I => \D_UU_AMIGA_in_6\
        );

    \I__1604\ : IoInMux
    port map (
            O => \N__6520\,
            I => \N__6517\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__6517\,
            I => \N__6514\
        );

    \I__1602\ : Span4Mux_s2_v
    port map (
            O => \N__6514\,
            I => \N__6511\
        );

    \I__1601\ : Span4Mux_h
    port map (
            O => \N__6511\,
            I => \N__6508\
        );

    \I__1600\ : Sp12to4
    port map (
            O => \N__6508\,
            I => \N__6505\
        );

    \I__1599\ : Span12Mux_s8_v
    port map (
            O => \N__6505\,
            I => \N__6502\
        );

    \I__1598\ : Odrv12
    port map (
            O => \N__6502\,
            I => \un1_D_UU_AMIGA_6\
        );

    \I__1597\ : IoInMux
    port map (
            O => \N__6499\,
            I => \N__6496\
        );

    \I__1596\ : LocalMux
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1595\ : Span4Mux_s2_h
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__1594\ : Sp12to4
    port map (
            O => \N__6490\,
            I => \N__6487\
        );

    \I__1593\ : Span12Mux_v
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__1592\ : Odrv12
    port map (
            O => \N__6484\,
            I => \un1_D_UM_AMIGA_2\
        );

    \I__1591\ : IoInMux
    port map (
            O => \N__6481\,
            I => \N__6478\
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__6478\,
            I => \N__6475\
        );

    \I__1589\ : Sp12to4
    port map (
            O => \N__6475\,
            I => \N__6472\
        );

    \I__1588\ : Span12Mux_h
    port map (
            O => \N__6472\,
            I => \N__6469\
        );

    \I__1587\ : Odrv12
    port map (
            O => \N__6469\,
            I => \un1_D_UM_AMIGA_6\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__6463\,
            I => \N__6460\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__6460\,
            I => \N__6455\
        );

    \I__1583\ : InMux
    port map (
            O => \N__6459\,
            I => \N__6452\
        );

    \I__1582\ : InMux
    port map (
            O => \N__6458\,
            I => \N__6449\
        );

    \I__1581\ : Span4Mux_v
    port map (
            O => \N__6455\,
            I => \N__6446\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__6452\,
            I => \N__6443\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__6449\,
            I => \N__6440\
        );

    \I__1578\ : Span4Mux_v
    port map (
            O => \N__6446\,
            I => \N__6433\
        );

    \I__1577\ : Span4Mux_v
    port map (
            O => \N__6443\,
            I => \N__6433\
        );

    \I__1576\ : Span4Mux_v
    port map (
            O => \N__6440\,
            I => \N__6433\
        );

    \I__1575\ : Sp12to4
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__1574\ : Span12Mux_h
    port map (
            O => \N__6430\,
            I => \N__6427\
        );

    \I__1573\ : Odrv12
    port map (
            O => \N__6427\,
            I => \D_UM_AMIGA_in_0\
        );

    \I__1572\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6421\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__6421\,
            I => \N__6418\
        );

    \I__1570\ : Odrv4
    port map (
            O => \N__6418\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\
        );

    \I__1569\ : InMux
    port map (
            O => \N__6415\,
            I => \N__6412\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N__6408\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6411\,
            I => \N__6405\
        );

    \I__1566\ : Span4Mux_v
    port map (
            O => \N__6408\,
            I => \N__6402\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6405\,
            I => \N__6398\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__6402\,
            I => \N__6395\
        );

    \I__1563\ : InMux
    port map (
            O => \N__6401\,
            I => \N__6392\
        );

    \I__1562\ : Span4Mux_v
    port map (
            O => \N__6398\,
            I => \N__6389\
        );

    \I__1561\ : Sp12to4
    port map (
            O => \N__6395\,
            I => \N__6382\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6392\,
            I => \N__6382\
        );

    \I__1559\ : Sp12to4
    port map (
            O => \N__6389\,
            I => \N__6382\
        );

    \I__1558\ : Span12Mux_h
    port map (
            O => \N__6382\,
            I => \N__6379\
        );

    \I__1557\ : Span12Mux_v
    port map (
            O => \N__6379\,
            I => \N__6376\
        );

    \I__1556\ : Odrv12
    port map (
            O => \N__6376\,
            I => \D_UM_AMIGA_in_6\
        );

    \I__1555\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6370\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__6370\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\
        );

    \I__1553\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__6361\,
            I => \N__6356\
        );

    \I__1550\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6353\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6350\
        );

    \I__1548\ : Span4Mux_v
    port map (
            O => \N__6356\,
            I => \N__6347\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__6353\,
            I => \N__6342\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6342\
        );

    \I__1545\ : Span4Mux_v
    port map (
            O => \N__6347\,
            I => \N__6339\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__6342\,
            I => \N__6336\
        );

    \I__1543\ : Sp12to4
    port map (
            O => \N__6339\,
            I => \N__6331\
        );

    \I__1542\ : Sp12to4
    port map (
            O => \N__6336\,
            I => \N__6331\
        );

    \I__1541\ : Span12Mux_h
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__6328\,
            I => \D_UM_AMIGA_in_2\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__1538\ : LocalMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__6319\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\
        );

    \I__1536\ : IoInMux
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6313\,
            I => \N__6310\
        );

    \I__1534\ : IoSpan4Mux
    port map (
            O => \N__6310\,
            I => \N__6307\
        );

    \I__1533\ : Span4Mux_s3_v
    port map (
            O => \N__6307\,
            I => \N__6304\
        );

    \I__1532\ : Span4Mux_v
    port map (
            O => \N__6304\,
            I => \N__6298\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6303\,
            I => \N__6295\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6302\,
            I => \N__6290\
        );

    \I__1529\ : InMux
    port map (
            O => \N__6301\,
            I => \N__6290\
        );

    \I__1528\ : Span4Mux_v
    port map (
            O => \N__6298\,
            I => \N__6283\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6295\,
            I => \N__6283\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6283\
        );

    \I__1525\ : Span4Mux_v
    port map (
            O => \N__6283\,
            I => \N__6279\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6282\,
            I => \N__6276\
        );

    \I__1523\ : Span4Mux_h
    port map (
            O => \N__6279\,
            I => \N__6272\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__6276\,
            I => \N__6269\
        );

    \I__1521\ : InMux
    port map (
            O => \N__6275\,
            I => \N__6266\
        );

    \I__1520\ : Sp12to4
    port map (
            O => \N__6272\,
            I => \N__6261\
        );

    \I__1519\ : Span12Mux_h
    port map (
            O => \N__6269\,
            I => \N__6261\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6258\
        );

    \I__1517\ : Span12Mux_v
    port map (
            O => \N__6261\,
            I => \N__6253\
        );

    \I__1516\ : Span12Mux_h
    port map (
            O => \N__6258\,
            I => \N__6253\
        );

    \I__1515\ : Odrv12
    port map (
            O => \N__6253\,
            I => \TACKn_in\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6250\,
            I => \N__6243\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6249\,
            I => \N__6236\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6248\,
            I => \N__6233\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6247\,
            I => \N__6228\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6246\,
            I => \N__6228\
        );

    \I__1509\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6225\
        );

    \I__1508\ : InMux
    port map (
            O => \N__6242\,
            I => \N__6218\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6241\,
            I => \N__6218\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6240\,
            I => \N__6218\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6215\
        );

    \I__1504\ : LocalMux
    port map (
            O => \N__6236\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6233\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6228\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__6225\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__6218\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6215\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__6202\,
            I => \N__6194\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6188\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6183\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6183\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6198\,
            I => \N__6178\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6197\,
            I => \N__6178\
        );

    \I__1492\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6175\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6170\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6170\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6167\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__6188\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6183\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6178\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6175\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6170\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__6167\,
            I => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__6154\,
            I => \N__6149\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6153\,
            I => \N__6144\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6141\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6138\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__6148\,
            I => \N__6134\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6147\,
            I => \N__6131\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6144\,
            I => \N__6122\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6141\,
            I => \N__6122\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__6138\,
            I => \N__6122\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6137\,
            I => \N__6117\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6117\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6131\,
            I => \N__6114\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6130\,
            I => \N__6109\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6129\,
            I => \N__6109\
        );

    \I__1468\ : Span4Mux_v
    port map (
            O => \N__6122\,
            I => \N__6106\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6117\,
            I => \N__6103\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__6114\,
            I => \N__6098\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__6109\,
            I => \N__6098\
        );

    \I__1464\ : Span4Mux_v
    port map (
            O => \N__6106\,
            I => \N__6095\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__6103\,
            I => \N__6089\
        );

    \I__1462\ : Span4Mux_v
    port map (
            O => \N__6098\,
            I => \N__6089\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__6095\,
            I => \N__6086\
        );

    \I__1460\ : InMux
    port map (
            O => \N__6094\,
            I => \N__6083\
        );

    \I__1459\ : Span4Mux_h
    port map (
            O => \N__6089\,
            I => \N__6080\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__6086\,
            I => \N__6075\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6075\
        );

    \I__1456\ : Sp12to4
    port map (
            O => \N__6080\,
            I => \N__6072\
        );

    \I__1455\ : Span4Mux_v
    port map (
            O => \N__6075\,
            I => \N__6069\
        );

    \I__1454\ : Span12Mux_s11_h
    port map (
            O => \N__6072\,
            I => \N__6066\
        );

    \I__1453\ : Span4Mux_h
    port map (
            O => \N__6069\,
            I => \N__6063\
        );

    \I__1452\ : Span12Mux_v
    port map (
            O => \N__6066\,
            I => \N__6058\
        );

    \I__1451\ : Sp12to4
    port map (
            O => \N__6063\,
            I => \N__6058\
        );

    \I__1450\ : Odrv12
    port map (
            O => \N__6058\,
            I => \RESETn_c\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__6055\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\
        );

    \I__1448\ : IoInMux
    port map (
            O => \N__6052\,
            I => \N__6049\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6049\,
            I => \N__6046\
        );

    \I__1446\ : Span4Mux_s3_v
    port map (
            O => \N__6046\,
            I => \N__6042\
        );

    \I__1445\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6038\
        );

    \I__1444\ : Span4Mux_h
    port map (
            O => \N__6042\,
            I => \N__6034\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6031\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6038\,
            I => \N__6028\
        );

    \I__1441\ : InMux
    port map (
            O => \N__6037\,
            I => \N__6025\
        );

    \I__1440\ : Span4Mux_v
    port map (
            O => \N__6034\,
            I => \N__6020\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6031\,
            I => \N__6020\
        );

    \I__1438\ : Span4Mux_h
    port map (
            O => \N__6028\,
            I => \N__6015\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6015\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__6020\,
            I => \N__6012\
        );

    \I__1435\ : Sp12to4
    port map (
            O => \N__6015\,
            I => \N__6009\
        );

    \I__1434\ : Sp12to4
    port map (
            O => \N__6012\,
            I => \N__6006\
        );

    \I__1433\ : Span12Mux_s11_v
    port map (
            O => \N__6009\,
            I => \N__6003\
        );

    \I__1432\ : Span12Mux_h
    port map (
            O => \N__6006\,
            I => \N__6000\
        );

    \I__1431\ : Span12Mux_h
    port map (
            O => \N__6003\,
            I => \N__5997\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__6000\,
            I => \RnW_c\
        );

    \I__1429\ : Odrv12
    port map (
            O => \N__5997\,
            I => \RnW_c\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__5992\,
            I => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_\
        );

    \I__1427\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5986\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__5986\,
            I => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\
        );

    \I__1425\ : InMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__5980\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\
        );

    \I__1423\ : InMux
    port map (
            O => \N__5977\,
            I => \N__5974\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__5974\,
            I => \N__5969\
        );

    \I__1421\ : InMux
    port map (
            O => \N__5973\,
            I => \N__5966\
        );

    \I__1420\ : InMux
    port map (
            O => \N__5972\,
            I => \N__5963\
        );

    \I__1419\ : Span4Mux_v
    port map (
            O => \N__5969\,
            I => \N__5960\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__5966\,
            I => \N__5955\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__5963\,
            I => \N__5955\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__5960\,
            I => \N__5952\
        );

    \I__1415\ : Span4Mux_v
    port map (
            O => \N__5955\,
            I => \N__5949\
        );

    \I__1414\ : Span4Mux_v
    port map (
            O => \N__5952\,
            I => \N__5946\
        );

    \I__1413\ : Span4Mux_v
    port map (
            O => \N__5949\,
            I => \N__5943\
        );

    \I__1412\ : Sp12to4
    port map (
            O => \N__5946\,
            I => \N__5938\
        );

    \I__1411\ : Sp12to4
    port map (
            O => \N__5943\,
            I => \N__5938\
        );

    \I__1410\ : Span12Mux_h
    port map (
            O => \N__5938\,
            I => \N__5935\
        );

    \I__1409\ : Odrv12
    port map (
            O => \N__5935\,
            I => \D_UU_AMIGA_in_1\
        );

    \I__1408\ : IoInMux
    port map (
            O => \N__5932\,
            I => \N__5929\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5926\
        );

    \I__1406\ : IoSpan4Mux
    port map (
            O => \N__5926\,
            I => \N__5923\
        );

    \I__1405\ : Span4Mux_s3_h
    port map (
            O => \N__5923\,
            I => \N__5920\
        );

    \I__1404\ : Sp12to4
    port map (
            O => \N__5920\,
            I => \N__5917\
        );

    \I__1403\ : Span12Mux_h
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__1402\ : Odrv12
    port map (
            O => \N__5914\,
            I => \un1_D_UU_AMIGA_1\
        );

    \I__1401\ : InMux
    port map (
            O => \N__5911\,
            I => \N__5908\
        );

    \I__1400\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5905\
        );

    \I__1399\ : Sp12to4
    port map (
            O => \N__5905\,
            I => \N__5900\
        );

    \I__1398\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5897\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__5903\,
            I => \N__5894\
        );

    \I__1396\ : Span12Mux_v
    port map (
            O => \N__5900\,
            I => \N__5891\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5888\
        );

    \I__1394\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5885\
        );

    \I__1393\ : Odrv12
    port map (
            O => \N__5891\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1392\ : Odrv4
    port map (
            O => \N__5888\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__5885\,
            I => \U111_CYCLE_SM.TA_ENZ0\
        );

    \I__1390\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__5875\,
            I => \N__5872\
        );

    \I__1388\ : Span4Mux_v
    port map (
            O => \N__5872\,
            I => \N__5868\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__5871\,
            I => \N__5863\
        );

    \I__1386\ : Span4Mux_v
    port map (
            O => \N__5868\,
            I => \N__5860\
        );

    \I__1385\ : InMux
    port map (
            O => \N__5867\,
            I => \N__5857\
        );

    \I__1384\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5854\
        );

    \I__1383\ : InMux
    port map (
            O => \N__5863\,
            I => \N__5851\
        );

    \I__1382\ : Span4Mux_v
    port map (
            O => \N__5860\,
            I => \N__5846\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__5857\,
            I => \N__5843\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__5854\,
            I => \N__5838\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__5851\,
            I => \N__5838\
        );

    \I__1378\ : InMux
    port map (
            O => \N__5850\,
            I => \N__5835\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__5849\,
            I => \N__5832\
        );

    \I__1376\ : Span4Mux_v
    port map (
            O => \N__5846\,
            I => \N__5828\
        );

    \I__1375\ : Span4Mux_v
    port map (
            O => \N__5843\,
            I => \N__5825\
        );

    \I__1374\ : Span4Mux_h
    port map (
            O => \N__5838\,
            I => \N__5822\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5819\
        );

    \I__1372\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5814\
        );

    \I__1371\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5814\
        );

    \I__1370\ : Sp12to4
    port map (
            O => \N__5828\,
            I => \N__5811\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__5825\,
            I => \N__5806\
        );

    \I__1368\ : Sp12to4
    port map (
            O => \N__5822\,
            I => \N__5806\
        );

    \I__1367\ : Span4Mux_h
    port map (
            O => \N__5819\,
            I => \N__5801\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5801\
        );

    \I__1365\ : Span12Mux_h
    port map (
            O => \N__5811\,
            I => \N__5796\
        );

    \I__1364\ : Span12Mux_v
    port map (
            O => \N__5806\,
            I => \N__5796\
        );

    \I__1363\ : Span4Mux_v
    port map (
            O => \N__5801\,
            I => \N__5793\
        );

    \I__1362\ : Odrv12
    port map (
            O => \N__5796\,
            I => \LBENn_c\
        );

    \I__1361\ : Odrv4
    port map (
            O => \N__5793\,
            I => \LBENn_c\
        );

    \I__1360\ : IoInMux
    port map (
            O => \N__5788\,
            I => \N__5785\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__1358\ : Span4Mux_s2_v
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__1357\ : Span4Mux_v
    port map (
            O => \N__5779\,
            I => \N__5776\
        );

    \I__1356\ : Span4Mux_v
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__5773\,
            I => \TAn_1_i\
        );

    \I__1354\ : InMux
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__5767\,
            I => \N__5763\
        );

    \I__1352\ : InMux
    port map (
            O => \N__5766\,
            I => \N__5760\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__5763\,
            I => \N__5757\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5754\
        );

    \I__1349\ : Sp12to4
    port map (
            O => \N__5757\,
            I => \N__5750\
        );

    \I__1348\ : Span4Mux_v
    port map (
            O => \N__5754\,
            I => \N__5747\
        );

    \I__1347\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5744\
        );

    \I__1346\ : Span12Mux_v
    port map (
            O => \N__5750\,
            I => \N__5741\
        );

    \I__1345\ : Sp12to4
    port map (
            O => \N__5747\,
            I => \N__5736\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5736\
        );

    \I__1343\ : Span12Mux_h
    port map (
            O => \N__5741\,
            I => \N__5733\
        );

    \I__1342\ : Span12Mux_h
    port map (
            O => \N__5736\,
            I => \N__5730\
        );

    \I__1341\ : Odrv12
    port map (
            O => \N__5733\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1340\ : Odrv12
    port map (
            O => \N__5730\,
            I => \D_UM_AMIGA_in_1\
        );

    \I__1339\ : InMux
    port map (
            O => \N__5725\,
            I => \N__5722\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__5722\,
            I => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\
        );

    \I__1337\ : IoInMux
    port map (
            O => \N__5719\,
            I => \N__5716\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__5716\,
            I => \N__5713\
        );

    \I__1335\ : Span4Mux_s3_h
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__1334\ : Sp12to4
    port map (
            O => \N__5710\,
            I => \N__5707\
        );

    \I__1333\ : Span12Mux_s10_v
    port map (
            O => \N__5707\,
            I => \N__5704\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__5704\,
            I => \un1_D_UM_AMIGA_1\
        );

    \I__1331\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5698\
        );

    \I__1330\ : LocalMux
    port map (
            O => \N__5698\,
            I => \N__5695\
        );

    \I__1329\ : Sp12to4
    port map (
            O => \N__5695\,
            I => \N__5692\
        );

    \I__1328\ : Odrv12
    port map (
            O => \N__5692\,
            I => \TS_CPUn_c\
        );

    \I__1327\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5683\
        );

    \I__1326\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5680\
        );

    \I__1325\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5677\
        );

    \I__1324\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5674\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__5683\,
            I => \N__5670\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5667\
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__5677\,
            I => \N__5664\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__5674\,
            I => \N__5661\
        );

    \I__1319\ : ClkMux
    port map (
            O => \N__5673\,
            I => \N__5650\
        );

    \I__1318\ : Glb2LocalMux
    port map (
            O => \N__5670\,
            I => \N__5650\
        );

    \I__1317\ : Glb2LocalMux
    port map (
            O => \N__5667\,
            I => \N__5650\
        );

    \I__1316\ : Glb2LocalMux
    port map (
            O => \N__5664\,
            I => \N__5650\
        );

    \I__1315\ : Glb2LocalMux
    port map (
            O => \N__5661\,
            I => \N__5650\
        );

    \I__1314\ : GlobalMux
    port map (
            O => \N__5650\,
            I => \CLK40\
        );

    \I__1313\ : InMux
    port map (
            O => \N__5647\,
            I => \N__5644\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__5644\,
            I => \N__5641\
        );

    \I__1311\ : Span4Mux_v
    port map (
            O => \N__5641\,
            I => \N__5638\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__5638\,
            I => \U111_CYCLE_SM.TS_EN_2_0\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5635\,
            I => \N__5632\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5632\,
            I => \N__5629\
        );

    \I__1307\ : Odrv12
    port map (
            O => \N__5629\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5626\,
            I => \N__5622\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5618\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5622\,
            I => \N__5615\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5621\,
            I => \N__5612\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5609\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__5615\,
            I => \N__5606\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__5612\,
            I => \N__5603\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__5609\,
            I => \N__5600\
        );

    \I__1298\ : Span4Mux_h
    port map (
            O => \N__5606\,
            I => \N__5597\
        );

    \I__1297\ : Span12Mux_h
    port map (
            O => \N__5603\,
            I => \N__5594\
        );

    \I__1296\ : Sp12to4
    port map (
            O => \N__5600\,
            I => \N__5589\
        );

    \I__1295\ : Sp12to4
    port map (
            O => \N__5597\,
            I => \N__5589\
        );

    \I__1294\ : Span12Mux_h
    port map (
            O => \N__5594\,
            I => \N__5586\
        );

    \I__1293\ : Span12Mux_h
    port map (
            O => \N__5589\,
            I => \N__5583\
        );

    \I__1292\ : Odrv12
    port map (
            O => \N__5586\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1291\ : Odrv12
    port map (
            O => \N__5583\,
            I => \D_UU_AMIGA_in_7\
        );

    \I__1290\ : IoInMux
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__1288\ : Span4Mux_s0_v
    port map (
            O => \N__5572\,
            I => \N__5569\
        );

    \I__1287\ : Span4Mux_v
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__5566\,
            I => \N__5563\
        );

    \I__1285\ : Sp12to4
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__1284\ : Odrv12
    port map (
            O => \N__5560\,
            I => \un1_D_UU_AMIGA_7\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5554\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__1281\ : Odrv12
    port map (
            O => \N__5551\,
            I => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\
        );

    \I__1280\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5544\
        );

    \I__1279\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5540\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5544\,
            I => \N__5537\
        );

    \I__1277\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5534\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__5540\,
            I => \N__5531\
        );

    \I__1275\ : Span4Mux_v
    port map (
            O => \N__5537\,
            I => \N__5528\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__5534\,
            I => \N__5525\
        );

    \I__1273\ : Sp12to4
    port map (
            O => \N__5531\,
            I => \N__5518\
        );

    \I__1272\ : Sp12to4
    port map (
            O => \N__5528\,
            I => \N__5518\
        );

    \I__1271\ : Span12Mux_s11_v
    port map (
            O => \N__5525\,
            I => \N__5518\
        );

    \I__1270\ : Span12Mux_h
    port map (
            O => \N__5518\,
            I => \N__5515\
        );

    \I__1269\ : Odrv12
    port map (
            O => \N__5515\,
            I => \D_UU_AMIGA_in_2\
        );

    \I__1268\ : IoInMux
    port map (
            O => \N__5512\,
            I => \N__5509\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5509\,
            I => \N__5506\
        );

    \I__1266\ : Span12Mux_s8_v
    port map (
            O => \N__5506\,
            I => \N__5503\
        );

    \I__1265\ : Odrv12
    port map (
            O => \N__5503\,
            I => \un1_D_UU_AMIGA_2\
        );

    \I__1264\ : IoInMux
    port map (
            O => \N__5500\,
            I => \N__5497\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__1262\ : IoSpan4Mux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__1261\ : Span4Mux_s3_h
    port map (
            O => \N__5491\,
            I => \N__5488\
        );

    \I__1260\ : Span4Mux_h
    port map (
            O => \N__5488\,
            I => \N__5485\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__5485\,
            I => \N__5482\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__5482\,
            I => \un1_D_UM_AMIGA_0\
        );

    \I__1257\ : InMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5473\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__1254\ : Span12Mux_v
    port map (
            O => \N__5470\,
            I => \N__5467\
        );

    \I__1253\ : Span12Mux_h
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__1252\ : Odrv12
    port map (
            O => \N__5464\,
            I => \BGn_c\
        );

    \I__1251\ : IoInMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5458\,
            I => \N__5453\
        );

    \I__1249\ : IoInMux
    port map (
            O => \N__5457\,
            I => \N__5449\
        );

    \I__1248\ : IoInMux
    port map (
            O => \N__5456\,
            I => \N__5446\
        );

    \I__1247\ : Span4Mux_s2_h
    port map (
            O => \N__5453\,
            I => \N__5443\
        );

    \I__1246\ : IoInMux
    port map (
            O => \N__5452\,
            I => \N__5440\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5430\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5446\,
            I => \N__5430\
        );

    \I__1243\ : IoSpan4Mux
    port map (
            O => \N__5443\,
            I => \N__5430\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__5440\,
            I => \N__5430\
        );

    \I__1241\ : IoInMux
    port map (
            O => \N__5439\,
            I => \N__5427\
        );

    \I__1240\ : IoSpan4Mux
    port map (
            O => \N__5430\,
            I => \N__5411\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5427\,
            I => \N__5411\
        );

    \I__1238\ : IoInMux
    port map (
            O => \N__5426\,
            I => \N__5408\
        );

    \I__1237\ : IoInMux
    port map (
            O => \N__5425\,
            I => \N__5405\
        );

    \I__1236\ : IoInMux
    port map (
            O => \N__5424\,
            I => \N__5402\
        );

    \I__1235\ : IoInMux
    port map (
            O => \N__5423\,
            I => \N__5399\
        );

    \I__1234\ : IoInMux
    port map (
            O => \N__5422\,
            I => \N__5396\
        );

    \I__1233\ : IoInMux
    port map (
            O => \N__5421\,
            I => \N__5393\
        );

    \I__1232\ : IoInMux
    port map (
            O => \N__5420\,
            I => \N__5389\
        );

    \I__1231\ : IoInMux
    port map (
            O => \N__5419\,
            I => \N__5386\
        );

    \I__1230\ : IoInMux
    port map (
            O => \N__5418\,
            I => \N__5378\
        );

    \I__1229\ : IoInMux
    port map (
            O => \N__5417\,
            I => \N__5375\
        );

    \I__1228\ : IoInMux
    port map (
            O => \N__5416\,
            I => \N__5372\
        );

    \I__1227\ : IoSpan4Mux
    port map (
            O => \N__5411\,
            I => \N__5357\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5357\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__5405\,
            I => \N__5357\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5357\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5399\,
            I => \N__5357\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5396\,
            I => \N__5357\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5393\,
            I => \N__5357\
        );

    \I__1220\ : IoInMux
    port map (
            O => \N__5392\,
            I => \N__5354\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5389\,
            I => \N__5347\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5347\
        );

    \I__1217\ : IoInMux
    port map (
            O => \N__5385\,
            I => \N__5344\
        );

    \I__1216\ : IoInMux
    port map (
            O => \N__5384\,
            I => \N__5341\
        );

    \I__1215\ : IoInMux
    port map (
            O => \N__5383\,
            I => \N__5338\
        );

    \I__1214\ : IoInMux
    port map (
            O => \N__5382\,
            I => \N__5335\
        );

    \I__1213\ : IoInMux
    port map (
            O => \N__5381\,
            I => \N__5332\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5378\,
            I => \N__5323\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5323\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5372\,
            I => \N__5323\
        );

    \I__1209\ : IoSpan4Mux
    port map (
            O => \N__5357\,
            I => \N__5317\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__5354\,
            I => \N__5317\
        );

    \I__1207\ : IoInMux
    port map (
            O => \N__5353\,
            I => \N__5314\
        );

    \I__1206\ : IoInMux
    port map (
            O => \N__5352\,
            I => \N__5310\
        );

    \I__1205\ : IoSpan4Mux
    port map (
            O => \N__5347\,
            I => \N__5299\
        );

    \I__1204\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5299\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__5341\,
            I => \N__5299\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5299\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__5335\,
            I => \N__5299\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__5332\,
            I => \N__5296\
        );

    \I__1199\ : IoInMux
    port map (
            O => \N__5331\,
            I => \N__5293\
        );

    \I__1198\ : IoInMux
    port map (
            O => \N__5330\,
            I => \N__5290\
        );

    \I__1197\ : IoSpan4Mux
    port map (
            O => \N__5323\,
            I => \N__5287\
        );

    \I__1196\ : IoInMux
    port map (
            O => \N__5322\,
            I => \N__5284\
        );

    \I__1195\ : IoSpan4Mux
    port map (
            O => \N__5317\,
            I => \N__5279\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5314\,
            I => \N__5279\
        );

    \I__1193\ : IoInMux
    port map (
            O => \N__5313\,
            I => \N__5276\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5310\,
            I => \N__5271\
        );

    \I__1191\ : IoSpan4Mux
    port map (
            O => \N__5299\,
            I => \N__5268\
        );

    \I__1190\ : Span4Mux_s3_v
    port map (
            O => \N__5296\,
            I => \N__5265\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5293\,
            I => \N__5259\
        );

    \I__1188\ : LocalMux
    port map (
            O => \N__5290\,
            I => \N__5259\
        );

    \I__1187\ : IoSpan4Mux
    port map (
            O => \N__5287\,
            I => \N__5254\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5284\,
            I => \N__5254\
        );

    \I__1185\ : IoSpan4Mux
    port map (
            O => \N__5279\,
            I => \N__5249\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5276\,
            I => \N__5249\
        );

    \I__1183\ : IoInMux
    port map (
            O => \N__5275\,
            I => \N__5246\
        );

    \I__1182\ : IoInMux
    port map (
            O => \N__5274\,
            I => \N__5243\
        );

    \I__1181\ : Span4Mux_s2_h
    port map (
            O => \N__5271\,
            I => \N__5236\
        );

    \I__1180\ : Span4Mux_s3_v
    port map (
            O => \N__5268\,
            I => \N__5236\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__5265\,
            I => \N__5236\
        );

    \I__1178\ : IoInMux
    port map (
            O => \N__5264\,
            I => \N__5233\
        );

    \I__1177\ : Span4Mux_s3_h
    port map (
            O => \N__5259\,
            I => \N__5230\
        );

    \I__1176\ : IoSpan4Mux
    port map (
            O => \N__5254\,
            I => \N__5225\
        );

    \I__1175\ : IoSpan4Mux
    port map (
            O => \N__5249\,
            I => \N__5225\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5246\,
            I => \N__5217\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5243\,
            I => \N__5217\
        );

    \I__1172\ : Sp12to4
    port map (
            O => \N__5236\,
            I => \N__5217\
        );

    \I__1171\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5214\
        );

    \I__1170\ : Span4Mux_v
    port map (
            O => \N__5230\,
            I => \N__5209\
        );

    \I__1169\ : Span4Mux_s3_h
    port map (
            O => \N__5225\,
            I => \N__5209\
        );

    \I__1168\ : IoInMux
    port map (
            O => \N__5224\,
            I => \N__5206\
        );

    \I__1167\ : Span12Mux_s11_v
    port map (
            O => \N__5217\,
            I => \N__5201\
        );

    \I__1166\ : Span12Mux_s2_h
    port map (
            O => \N__5214\,
            I => \N__5201\
        );

    \I__1165\ : Sp12to4
    port map (
            O => \N__5209\,
            I => \N__5196\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5196\
        );

    \I__1163\ : Span12Mux_h
    port map (
            O => \N__5201\,
            I => \N__5193\
        );

    \I__1162\ : Span12Mux_s8_h
    port map (
            O => \N__5196\,
            I => \N__5190\
        );

    \I__1161\ : Odrv12
    port map (
            O => \N__5193\,
            I => \CPU_READ_EN_i\
        );

    \I__1160\ : Odrv12
    port map (
            O => \N__5190\,
            I => \CPU_READ_EN_i\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__5185\,
            I => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\
        );

    \I__1158\ : CascadeMux
    port map (
            O => \N__5182\,
            I => \N__5177\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5172\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5180\,
            I => \N__5167\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5177\,
            I => \N__5167\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5162\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5162\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5172\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__5167\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5162\,
            I => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\
        );

    \I__1149\ : CascadeMux
    port map (
            O => \N__5155\,
            I => \U111_CYCLE_SM.N_97_cascade_\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5152\,
            I => \N__5149\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__5149\,
            I => \U111_CYCLE_SM.LW_CYCLE_0\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5146\,
            I => \N__5143\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__1144\ : Span12Mux_h
    port map (
            O => \N__5140\,
            I => \N__5135\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5139\,
            I => \N__5130\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5130\
        );

    \I__1141\ : Span12Mux_v
    port map (
            O => \N__5135\,
            I => \N__5127\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5130\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__1139\ : Odrv12
    port map (
            O => \N__5127\,
            I => \U111_CYCLE_SM.TS_ENZ0\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5119\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5119\,
            I => \U111_CYCLE_SM.un3_LW_CYCLE_START\
        );

    \I__1136\ : SRMux
    port map (
            O => \N__5116\,
            I => \N__5113\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__1134\ : Span4Mux_h
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__1133\ : Odrv4
    port map (
            O => \N__5107\,
            I => \U111_CYCLE_SM.RESETn_c_i\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5104\,
            I => \N__5101\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5101\,
            I => \N__5098\
        );

    \I__1130\ : Span4Mux_v
    port map (
            O => \N__5098\,
            I => \N__5095\
        );

    \I__1129\ : Sp12to4
    port map (
            O => \N__5095\,
            I => \N__5092\
        );

    \I__1128\ : Span12Mux_h
    port map (
            O => \N__5092\,
            I => \N__5089\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__5089\,
            I => \SIZ_c_1\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5083\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__1124\ : Span4Mux_v
    port map (
            O => \N__5080\,
            I => \N__5077\
        );

    \I__1123\ : Sp12to4
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__1122\ : Span12Mux_h
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__1121\ : Odrv12
    port map (
            O => \N__5071\,
            I => \SIZ_c_0\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5068\,
            I => \N__5065\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5061\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5064\,
            I => \N__5058\
        );

    \I__1117\ : Span4Mux_v
    port map (
            O => \N__5061\,
            I => \N__5053\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__5058\,
            I => \N__5053\
        );

    \I__1115\ : Span4Mux_v
    port map (
            O => \N__5053\,
            I => \N__5050\
        );

    \I__1114\ : Sp12to4
    port map (
            O => \N__5050\,
            I => \N__5047\
        );

    \I__1113\ : Span12Mux_h
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__1112\ : Span12Mux_v
    port map (
            O => \N__5044\,
            I => \N__5041\
        );

    \I__1111\ : Odrv12
    port map (
            O => \N__5041\,
            I => \PORTSIZE_c\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5034\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5031\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5034\,
            I => \N__5028\
        );

    \I__1107\ : LocalMux
    port map (
            O => \N__5031\,
            I => \N__5025\
        );

    \I__1106\ : Odrv12
    port map (
            O => \N__5028\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1105\ : Odrv12
    port map (
            O => \N__5025\,
            I => \U111_CYCLE_SM.LW_TRANS_0\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5020\,
            I => \N__5017\
        );

    \I__1103\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__5014\
        );

    \I__1102\ : Span4Mux_v
    port map (
            O => \N__5014\,
            I => \N__5011\
        );

    \I__1101\ : Sp12to4
    port map (
            O => \N__5011\,
            I => \N__5008\
        );

    \I__1100\ : Span12Mux_h
    port map (
            O => \N__5008\,
            I => \N__5005\
        );

    \I__1099\ : Odrv12
    port map (
            O => \N__5005\,
            I => \D_LM_AMIGA_in_7\
        );

    \I__1098\ : IoInMux
    port map (
            O => \N__5002\,
            I => \N__4999\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__4999\,
            I => \N__4996\
        );

    \I__1096\ : IoSpan4Mux
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__1095\ : Span4Mux_s2_h
    port map (
            O => \N__4993\,
            I => \N__4990\
        );

    \I__1094\ : Sp12to4
    port map (
            O => \N__4990\,
            I => \N__4987\
        );

    \I__1093\ : Odrv12
    port map (
            O => \N__4987\,
            I => \un1_D_LM_AMIGA_7\
        );

    \I__1092\ : IoInMux
    port map (
            O => \N__4984\,
            I => \N__4981\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__4981\,
            I => \N__4977\
        );

    \I__1090\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4974\
        );

    \I__1089\ : IoSpan4Mux
    port map (
            O => \N__4977\,
            I => \N__4971\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__4974\,
            I => \N__4968\
        );

    \I__1087\ : Span4Mux_s3_h
    port map (
            O => \N__4971\,
            I => \N__4965\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__4968\,
            I => \N__4962\
        );

    \I__1085\ : Sp12to4
    port map (
            O => \N__4965\,
            I => \N__4959\
        );

    \I__1084\ : Sp12to4
    port map (
            O => \N__4962\,
            I => \N__4956\
        );

    \I__1083\ : Span12Mux_v
    port map (
            O => \N__4959\,
            I => \N__4953\
        );

    \I__1082\ : Span12Mux_v
    port map (
            O => \N__4956\,
            I => \N__4950\
        );

    \I__1081\ : Span12Mux_h
    port map (
            O => \N__4953\,
            I => \N__4947\
        );

    \I__1080\ : Span12Mux_v
    port map (
            O => \N__4950\,
            I => \N__4944\
        );

    \I__1079\ : Span12Mux_h
    port map (
            O => \N__4947\,
            I => \N__4941\
        );

    \I__1078\ : Span12Mux_h
    port map (
            O => \N__4944\,
            I => \N__4938\
        );

    \I__1077\ : Odrv12
    port map (
            O => \N__4941\,
            I => \D_LL_040_in_5\
        );

    \I__1076\ : Odrv12
    port map (
            O => \N__4938\,
            I => \D_LL_040_in_5\
        );

    \I__1075\ : InMux
    port map (
            O => \N__4933\,
            I => \N__4930\
        );

    \I__1074\ : LocalMux
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__4927\,
            I => \N__4924\
        );

    \I__1072\ : Sp12to4
    port map (
            O => \N__4924\,
            I => \N__4921\
        );

    \I__1071\ : Span12Mux_h
    port map (
            O => \N__4921\,
            I => \N__4918\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__4918\,
            I => \D_UM_040_in_5\
        );

    \I__1069\ : IoInMux
    port map (
            O => \N__4915\,
            I => \N__4912\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__4912\,
            I => \N__4909\
        );

    \I__1067\ : Span12Mux_s10_v
    port map (
            O => \N__4909\,
            I => \N__4906\
        );

    \I__1066\ : Span12Mux_h
    port map (
            O => \N__4906\,
            I => \N__4903\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__4903\,
            I => \un1_D_UM_040_5\
        );

    \I__1064\ : InMux
    port map (
            O => \N__4900\,
            I => \N__4897\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__4897\,
            I => \N__4894\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__1061\ : Sp12to4
    port map (
            O => \N__4891\,
            I => \N__4888\
        );

    \I__1060\ : Span12Mux_h
    port map (
            O => \N__4888\,
            I => \N__4885\
        );

    \I__1059\ : Odrv12
    port map (
            O => \N__4885\,
            I => \D_UU_040_in_3\
        );

    \I__1058\ : InMux
    port map (
            O => \N__4882\,
            I => \N__4875\
        );

    \I__1057\ : InMux
    port map (
            O => \N__4881\,
            I => \N__4872\
        );

    \I__1056\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4864\
        );

    \I__1055\ : InMux
    port map (
            O => \N__4879\,
            I => \N__4864\
        );

    \I__1054\ : InMux
    port map (
            O => \N__4878\,
            I => \N__4861\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__4875\,
            I => \N__4850\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__4872\,
            I => \N__4850\
        );

    \I__1051\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4847\
        );

    \I__1050\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4844\
        );

    \I__1049\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4841\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__4864\,
            I => \N__4836\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__4861\,
            I => \N__4836\
        );

    \I__1046\ : InMux
    port map (
            O => \N__4860\,
            I => \N__4831\
        );

    \I__1045\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4831\
        );

    \I__1044\ : InMux
    port map (
            O => \N__4858\,
            I => \N__4824\
        );

    \I__1043\ : InMux
    port map (
            O => \N__4857\,
            I => \N__4824\
        );

    \I__1042\ : InMux
    port map (
            O => \N__4856\,
            I => \N__4821\
        );

    \I__1041\ : InMux
    port map (
            O => \N__4855\,
            I => \N__4809\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__4850\,
            I => \N__4800\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__4847\,
            I => \N__4800\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__4844\,
            I => \N__4800\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4797\
        );

    \I__1036\ : Span4Mux_v
    port map (
            O => \N__4836\,
            I => \N__4792\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__4831\,
            I => \N__4792\
        );

    \I__1034\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4789\
        );

    \I__1033\ : InMux
    port map (
            O => \N__4829\,
            I => \N__4786\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__4824\,
            I => \N__4781\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__4821\,
            I => \N__4781\
        );

    \I__1030\ : InMux
    port map (
            O => \N__4820\,
            I => \N__4778\
        );

    \I__1029\ : InMux
    port map (
            O => \N__4819\,
            I => \N__4775\
        );

    \I__1028\ : InMux
    port map (
            O => \N__4818\,
            I => \N__4770\
        );

    \I__1027\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4770\
        );

    \I__1026\ : InMux
    port map (
            O => \N__4816\,
            I => \N__4765\
        );

    \I__1025\ : InMux
    port map (
            O => \N__4815\,
            I => \N__4765\
        );

    \I__1024\ : InMux
    port map (
            O => \N__4814\,
            I => \N__4762\
        );

    \I__1023\ : InMux
    port map (
            O => \N__4813\,
            I => \N__4754\
        );

    \I__1022\ : InMux
    port map (
            O => \N__4812\,
            I => \N__4754\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__4809\,
            I => \N__4751\
        );

    \I__1020\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4746\
        );

    \I__1019\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4746\
        );

    \I__1018\ : Span4Mux_v
    port map (
            O => \N__4800\,
            I => \N__4743\
        );

    \I__1017\ : Span4Mux_v
    port map (
            O => \N__4797\,
            I => \N__4734\
        );

    \I__1016\ : Span4Mux_v
    port map (
            O => \N__4792\,
            I => \N__4734\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__4789\,
            I => \N__4734\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__4786\,
            I => \N__4734\
        );

    \I__1013\ : Span4Mux_v
    port map (
            O => \N__4781\,
            I => \N__4729\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__4778\,
            I => \N__4729\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__4775\,
            I => \N__4726\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__4770\,
            I => \N__4723\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__4765\,
            I => \N__4720\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__4762\,
            I => \N__4717\
        );

    \I__1007\ : InMux
    port map (
            O => \N__4761\,
            I => \N__4712\
        );

    \I__1006\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4712\
        );

    \I__1005\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4709\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__4754\,
            I => \N__4705\
        );

    \I__1003\ : Span12Mux_h
    port map (
            O => \N__4751\,
            I => \N__4700\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__4746\,
            I => \N__4700\
        );

    \I__1001\ : Span4Mux_v
    port map (
            O => \N__4743\,
            I => \N__4697\
        );

    \I__1000\ : Span4Mux_v
    port map (
            O => \N__4734\,
            I => \N__4694\
        );

    \I__999\ : Span4Mux_v
    port map (
            O => \N__4729\,
            I => \N__4687\
        );

    \I__998\ : Span4Mux_v
    port map (
            O => \N__4726\,
            I => \N__4687\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__4723\,
            I => \N__4687\
        );

    \I__996\ : Span4Mux_v
    port map (
            O => \N__4720\,
            I => \N__4680\
        );

    \I__995\ : Span4Mux_h
    port map (
            O => \N__4717\,
            I => \N__4680\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__4712\,
            I => \N__4680\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__4709\,
            I => \N__4677\
        );

    \I__992\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4674\
        );

    \I__991\ : Odrv12
    port map (
            O => \N__4705\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__990\ : Odrv12
    port map (
            O => \N__4700\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__989\ : Odrv4
    port map (
            O => \N__4697\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__988\ : Odrv4
    port map (
            O => \N__4694\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__4687\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__4680\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__985\ : Odrv12
    port map (
            O => \N__4677\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__4674\,
            I => \U111_CYCLE_SM.FLIP\
        );

    \I__983\ : IoInMux
    port map (
            O => \N__4657\,
            I => \N__4654\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__4654\,
            I => \N__4651\
        );

    \I__981\ : IoSpan4Mux
    port map (
            O => \N__4651\,
            I => \N__4647\
        );

    \I__980\ : InMux
    port map (
            O => \N__4650\,
            I => \N__4644\
        );

    \I__979\ : IoSpan4Mux
    port map (
            O => \N__4647\,
            I => \N__4641\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__4644\,
            I => \N__4638\
        );

    \I__977\ : Span4Mux_s2_h
    port map (
            O => \N__4641\,
            I => \N__4635\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__4638\,
            I => \N__4632\
        );

    \I__975\ : Sp12to4
    port map (
            O => \N__4635\,
            I => \N__4629\
        );

    \I__974\ : Sp12to4
    port map (
            O => \N__4632\,
            I => \N__4626\
        );

    \I__973\ : Span12Mux_h
    port map (
            O => \N__4629\,
            I => \N__4623\
        );

    \I__972\ : Span12Mux_v
    port map (
            O => \N__4626\,
            I => \N__4620\
        );

    \I__971\ : Span12Mux_h
    port map (
            O => \N__4623\,
            I => \N__4617\
        );

    \I__970\ : Span12Mux_h
    port map (
            O => \N__4620\,
            I => \N__4614\
        );

    \I__969\ : Odrv12
    port map (
            O => \N__4617\,
            I => \D_LM_040_in_3\
        );

    \I__968\ : Odrv12
    port map (
            O => \N__4614\,
            I => \D_LM_040_in_3\
        );

    \I__967\ : IoInMux
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__4606\,
            I => \N__4603\
        );

    \I__965\ : IoSpan4Mux
    port map (
            O => \N__4603\,
            I => \N__4600\
        );

    \I__964\ : IoSpan4Mux
    port map (
            O => \N__4600\,
            I => \N__4597\
        );

    \I__963\ : Span4Mux_s2_v
    port map (
            O => \N__4597\,
            I => \N__4594\
        );

    \I__962\ : Span4Mux_h
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__961\ : Span4Mux_v
    port map (
            O => \N__4591\,
            I => \N__4588\
        );

    \I__960\ : Odrv4
    port map (
            O => \N__4588\,
            I => \un1_D_UU_040_3\
        );

    \I__959\ : IoInMux
    port map (
            O => \N__4585\,
            I => \N__4582\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4582\,
            I => \N__4579\
        );

    \I__957\ : Span4Mux_s2_v
    port map (
            O => \N__4579\,
            I => \N__4576\
        );

    \I__956\ : Span4Mux_v
    port map (
            O => \N__4576\,
            I => \N__4573\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__4573\,
            I => \N__4570\
        );

    \I__954\ : Span4Mux_h
    port map (
            O => \N__4570\,
            I => \N__4567\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__4567\,
            I => \U111_CYCLE_SM_TBI_CPUn_0_i\
        );

    \I__952\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4561\,
            I => \U111_CYCLE_SM.TS_EN_5\
        );

    \I__950\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__4555\,
            I => \N__4552\
        );

    \I__948\ : Span12Mux_h
    port map (
            O => \N__4552\,
            I => \N__4549\
        );

    \I__947\ : Odrv12
    port map (
            O => \N__4549\,
            I => \D_LM_AMIGA_in_1\
        );

    \I__946\ : CascadeMux
    port map (
            O => \N__4546\,
            I => \U111_CYCLE_SM.FLIP_cascade_\
        );

    \I__945\ : IoInMux
    port map (
            O => \N__4543\,
            I => \N__4540\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__943\ : Span4Mux_s3_h
    port map (
            O => \N__4537\,
            I => \N__4534\
        );

    \I__942\ : Sp12to4
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__941\ : Span12Mux_v
    port map (
            O => \N__4531\,
            I => \N__4528\
        );

    \I__940\ : Odrv12
    port map (
            O => \N__4528\,
            I => \un1_D_LM_AMIGA_1\
        );

    \I__939\ : IoInMux
    port map (
            O => \N__4525\,
            I => \N__4522\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__937\ : IoInMux
    port map (
            O => \N__4521\,
            I => \N__4513\
        );

    \I__936\ : IoInMux
    port map (
            O => \N__4520\,
            I => \N__4510\
        );

    \I__935\ : IoInMux
    port map (
            O => \N__4519\,
            I => \N__4507\
        );

    \I__934\ : IoSpan4Mux
    port map (
            O => \N__4516\,
            I => \N__4504\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4513\,
            I => \N__4501\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__4510\,
            I => \N__4498\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4507\,
            I => \N__4495\
        );

    \I__930\ : IoSpan4Mux
    port map (
            O => \N__4504\,
            I => \N__4490\
        );

    \I__929\ : IoSpan4Mux
    port map (
            O => \N__4501\,
            I => \N__4490\
        );

    \I__928\ : IoSpan4Mux
    port map (
            O => \N__4498\,
            I => \N__4487\
        );

    \I__927\ : IoSpan4Mux
    port map (
            O => \N__4495\,
            I => \N__4484\
        );

    \I__926\ : Span4Mux_s2_v
    port map (
            O => \N__4490\,
            I => \N__4481\
        );

    \I__925\ : Sp12to4
    port map (
            O => \N__4487\,
            I => \N__4478\
        );

    \I__924\ : Sp12to4
    port map (
            O => \N__4484\,
            I => \N__4475\
        );

    \I__923\ : Sp12to4
    port map (
            O => \N__4481\,
            I => \N__4472\
        );

    \I__922\ : Span12Mux_h
    port map (
            O => \N__4478\,
            I => \N__4467\
        );

    \I__921\ : Span12Mux_s7_h
    port map (
            O => \N__4475\,
            I => \N__4467\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__4472\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__919\ : Odrv12
    port map (
            O => \N__4467\,
            I => \GB_BUFFER_CLK40_THRU_CO\
        );

    \I__918\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4459\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__4459\,
            I => \N__4455\
        );

    \I__916\ : ClkMux
    port map (
            O => \N__4458\,
            I => \N__4429\
        );

    \I__915\ : Glb2LocalMux
    port map (
            O => \N__4455\,
            I => \N__4429\
        );

    \I__914\ : ClkMux
    port map (
            O => \N__4454\,
            I => \N__4429\
        );

    \I__913\ : ClkMux
    port map (
            O => \N__4453\,
            I => \N__4429\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4452\,
            I => \N__4429\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4451\,
            I => \N__4429\
        );

    \I__910\ : ClkMux
    port map (
            O => \N__4450\,
            I => \N__4429\
        );

    \I__909\ : ClkMux
    port map (
            O => \N__4449\,
            I => \N__4429\
        );

    \I__908\ : ClkMux
    port map (
            O => \N__4448\,
            I => \N__4429\
        );

    \I__907\ : GlobalMux
    port map (
            O => \N__4429\,
            I => \CLK80\
        );

    \I__906\ : IoInMux
    port map (
            O => \N__4426\,
            I => \N__4423\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__4423\,
            I => \N__4419\
        );

    \I__904\ : IoInMux
    port map (
            O => \N__4422\,
            I => \N__4416\
        );

    \I__903\ : Span12Mux_s2_v
    port map (
            O => \N__4419\,
            I => \N__4413\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__4416\,
            I => \N__4410\
        );

    \I__901\ : Span12Mux_v
    port map (
            O => \N__4413\,
            I => \N__4407\
        );

    \I__900\ : Span12Mux_s9_h
    port map (
            O => \N__4410\,
            I => \N__4404\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__4407\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__898\ : Odrv12
    port map (
            O => \N__4404\,
            I => \GB_BUFFER_CLK80_THRU_CO\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__4399\,
            I => \U111_CYCLE_SM.A_OUT_0_cascade_\
        );

    \I__896\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4393\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4393\,
            I => \N__4390\
        );

    \I__894\ : Span12Mux_s10_h
    port map (
            O => \N__4390\,
            I => \N__4387\
        );

    \I__893\ : Span12Mux_v
    port map (
            O => \N__4387\,
            I => \N__4383\
        );

    \I__892\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4380\
        );

    \I__891\ : Odrv12
    port map (
            O => \N__4383\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__4380\,
            I => \U111_CYCLE_SM.A_OUTZ0\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__4375\,
            I => \U111_CYCLE_SM.N_75_0_cascade_\
        );

    \I__888\ : IoInMux
    port map (
            O => \N__4372\,
            I => \N__4369\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__4369\,
            I => \N__4366\
        );

    \I__886\ : Span4Mux_s3_h
    port map (
            O => \N__4366\,
            I => \N__4363\
        );

    \I__885\ : Span4Mux_v
    port map (
            O => \N__4363\,
            I => \N__4360\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__4360\,
            I => \N__4357\
        );

    \I__883\ : Span12Mux_h
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__4354\,
            I => \un1_D_LM_AMIGA_0\
        );

    \I__881\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4348\,
            I => \N__4345\
        );

    \I__879\ : Span12Mux_v
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__878\ : Span12Mux_h
    port map (
            O => \N__4342\,
            I => \N__4339\
        );

    \I__877\ : Odrv12
    port map (
            O => \N__4339\,
            I => \D_LL_AMIGA_in_7\
        );

    \I__876\ : IoInMux
    port map (
            O => \N__4336\,
            I => \N__4333\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4333\,
            I => \N__4330\
        );

    \I__874\ : Span4Mux_s3_h
    port map (
            O => \N__4330\,
            I => \N__4327\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__4327\,
            I => \N__4324\
        );

    \I__872\ : Span4Mux_v
    port map (
            O => \N__4324\,
            I => \N__4321\
        );

    \I__871\ : Sp12to4
    port map (
            O => \N__4321\,
            I => \N__4318\
        );

    \I__870\ : Odrv12
    port map (
            O => \N__4318\,
            I => \un1_D_LL_AMIGA_7\
        );

    \I__869\ : IoInMux
    port map (
            O => \N__4315\,
            I => \N__4312\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4312\,
            I => \N__4308\
        );

    \I__867\ : InMux
    port map (
            O => \N__4311\,
            I => \N__4305\
        );

    \I__866\ : IoSpan4Mux
    port map (
            O => \N__4308\,
            I => \N__4302\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4299\
        );

    \I__864\ : Span4Mux_s2_h
    port map (
            O => \N__4302\,
            I => \N__4296\
        );

    \I__863\ : Span4Mux_v
    port map (
            O => \N__4299\,
            I => \N__4293\
        );

    \I__862\ : Sp12to4
    port map (
            O => \N__4296\,
            I => \N__4290\
        );

    \I__861\ : Sp12to4
    port map (
            O => \N__4293\,
            I => \N__4287\
        );

    \I__860\ : Span12Mux_h
    port map (
            O => \N__4290\,
            I => \N__4284\
        );

    \I__859\ : Span12Mux_h
    port map (
            O => \N__4287\,
            I => \N__4281\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__4284\,
            I => \N__4278\
        );

    \I__857\ : Span12Mux_v
    port map (
            O => \N__4281\,
            I => \N__4275\
        );

    \I__856\ : Odrv12
    port map (
            O => \N__4278\,
            I => \D_LL_040_in_0\
        );

    \I__855\ : Odrv12
    port map (
            O => \N__4275\,
            I => \D_LL_040_in_0\
        );

    \I__854\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__4267\,
            I => \N__4264\
        );

    \I__852\ : Span12Mux_h
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__851\ : Odrv12
    port map (
            O => \N__4261\,
            I => \D_UM_040_in_0\
        );

    \I__850\ : IoInMux
    port map (
            O => \N__4258\,
            I => \N__4255\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__4255\,
            I => \N__4252\
        );

    \I__848\ : IoSpan4Mux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__847\ : Span4Mux_s0_h
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__846\ : Sp12to4
    port map (
            O => \N__4246\,
            I => \N__4243\
        );

    \I__845\ : Span12Mux_s11_h
    port map (
            O => \N__4243\,
            I => \N__4240\
        );

    \I__844\ : Odrv12
    port map (
            O => \N__4240\,
            I => \un1_D_UM_040_0\
        );

    \I__843\ : InMux
    port map (
            O => \N__4237\,
            I => \N__4234\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4231\
        );

    \I__841\ : Span4Mux_h
    port map (
            O => \N__4231\,
            I => \N__4228\
        );

    \I__840\ : Sp12to4
    port map (
            O => \N__4228\,
            I => \N__4225\
        );

    \I__839\ : Span12Mux_v
    port map (
            O => \N__4225\,
            I => \N__4222\
        );

    \I__838\ : Span12Mux_h
    port map (
            O => \N__4222\,
            I => \N__4219\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__4219\,
            I => \D_UM_040_in_4\
        );

    \I__836\ : InMux
    port map (
            O => \N__4216\,
            I => \N__4212\
        );

    \I__835\ : IoInMux
    port map (
            O => \N__4215\,
            I => \N__4209\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__4212\,
            I => \N__4206\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__4209\,
            I => \N__4203\
        );

    \I__832\ : Span4Mux_v
    port map (
            O => \N__4206\,
            I => \N__4200\
        );

    \I__831\ : Span4Mux_s2_h
    port map (
            O => \N__4203\,
            I => \N__4197\
        );

    \I__830\ : Sp12to4
    port map (
            O => \N__4200\,
            I => \N__4194\
        );

    \I__829\ : Span4Mux_v
    port map (
            O => \N__4197\,
            I => \N__4191\
        );

    \I__828\ : Span12Mux_h
    port map (
            O => \N__4194\,
            I => \N__4188\
        );

    \I__827\ : Sp12to4
    port map (
            O => \N__4191\,
            I => \N__4185\
        );

    \I__826\ : Span12Mux_v
    port map (
            O => \N__4188\,
            I => \N__4182\
        );

    \I__825\ : Span12Mux_h
    port map (
            O => \N__4185\,
            I => \N__4179\
        );

    \I__824\ : Span12Mux_v
    port map (
            O => \N__4182\,
            I => \N__4176\
        );

    \I__823\ : Span12Mux_h
    port map (
            O => \N__4179\,
            I => \N__4173\
        );

    \I__822\ : Odrv12
    port map (
            O => \N__4176\,
            I => \D_LL_040_in_4\
        );

    \I__821\ : Odrv12
    port map (
            O => \N__4173\,
            I => \D_LL_040_in_4\
        );

    \I__820\ : IoInMux
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4165\,
            I => \N__4162\
        );

    \I__818\ : Span12Mux_s3_h
    port map (
            O => \N__4162\,
            I => \N__4159\
        );

    \I__817\ : Span12Mux_h
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__4156\,
            I => \un1_D_UM_040_4\
        );

    \I__815\ : IoInMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__4150\,
            I => \N__4147\
        );

    \I__813\ : IoSpan4Mux
    port map (
            O => \N__4147\,
            I => \N__4143\
        );

    \I__812\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4140\
        );

    \I__811\ : Span4Mux_s0_h
    port map (
            O => \N__4143\,
            I => \N__4137\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4140\,
            I => \N__4134\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__4137\,
            I => \N__4131\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__4134\,
            I => \N__4128\
        );

    \I__807\ : Sp12to4
    port map (
            O => \N__4131\,
            I => \N__4125\
        );

    \I__806\ : Sp12to4
    port map (
            O => \N__4128\,
            I => \N__4122\
        );

    \I__805\ : Span12Mux_h
    port map (
            O => \N__4125\,
            I => \N__4119\
        );

    \I__804\ : Span12Mux_h
    port map (
            O => \N__4122\,
            I => \N__4116\
        );

    \I__803\ : Span12Mux_h
    port map (
            O => \N__4119\,
            I => \N__4113\
        );

    \I__802\ : Span12Mux_v
    port map (
            O => \N__4116\,
            I => \N__4110\
        );

    \I__801\ : Odrv12
    port map (
            O => \N__4113\,
            I => \D_LM_040_in_5\
        );

    \I__800\ : Odrv12
    port map (
            O => \N__4110\,
            I => \D_LM_040_in_5\
        );

    \I__799\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4102\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4102\,
            I => \N__4099\
        );

    \I__797\ : Span4Mux_v
    port map (
            O => \N__4099\,
            I => \N__4096\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__4096\,
            I => \N__4093\
        );

    \I__795\ : Sp12to4
    port map (
            O => \N__4093\,
            I => \N__4090\
        );

    \I__794\ : Span12Mux_h
    port map (
            O => \N__4090\,
            I => \N__4087\
        );

    \I__793\ : Odrv12
    port map (
            O => \N__4087\,
            I => \D_UU_040_in_5\
        );

    \I__792\ : IoInMux
    port map (
            O => \N__4084\,
            I => \N__4081\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4081\,
            I => \N__4078\
        );

    \I__790\ : Span4Mux_s3_h
    port map (
            O => \N__4078\,
            I => \N__4075\
        );

    \I__789\ : Sp12to4
    port map (
            O => \N__4075\,
            I => \N__4072\
        );

    \I__788\ : Span12Mux_s10_v
    port map (
            O => \N__4072\,
            I => \N__4069\
        );

    \I__787\ : Span12Mux_h
    port map (
            O => \N__4069\,
            I => \N__4066\
        );

    \I__786\ : Odrv12
    port map (
            O => \N__4066\,
            I => \un1_D_UU_040_5\
        );

    \I__785\ : IoInMux
    port map (
            O => \N__4063\,
            I => \N__4060\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__4060\,
            I => \N__4057\
        );

    \I__783\ : IoSpan4Mux
    port map (
            O => \N__4057\,
            I => \N__4053\
        );

    \I__782\ : InMux
    port map (
            O => \N__4056\,
            I => \N__4050\
        );

    \I__781\ : Span4Mux_s2_h
    port map (
            O => \N__4053\,
            I => \N__4047\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4050\,
            I => \N__4044\
        );

    \I__779\ : Sp12to4
    port map (
            O => \N__4047\,
            I => \N__4041\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__4044\,
            I => \N__4038\
        );

    \I__777\ : Span12Mux_h
    port map (
            O => \N__4041\,
            I => \N__4035\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__4038\,
            I => \N__4032\
        );

    \I__775\ : Span12Mux_h
    port map (
            O => \N__4035\,
            I => \N__4029\
        );

    \I__774\ : Sp12to4
    port map (
            O => \N__4032\,
            I => \N__4026\
        );

    \I__773\ : Odrv12
    port map (
            O => \N__4029\,
            I => \D_LM_040_in_7\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__4026\,
            I => \D_LM_040_in_7\
        );

    \I__771\ : InMux
    port map (
            O => \N__4021\,
            I => \N__4018\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4018\,
            I => \N__4015\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__4015\,
            I => \N__4012\
        );

    \I__768\ : Sp12to4
    port map (
            O => \N__4012\,
            I => \N__4009\
        );

    \I__767\ : Span12Mux_h
    port map (
            O => \N__4009\,
            I => \N__4006\
        );

    \I__766\ : Odrv12
    port map (
            O => \N__4006\,
            I => \D_UU_040_in_7\
        );

    \I__765\ : IoInMux
    port map (
            O => \N__4003\,
            I => \N__4000\
        );

    \I__764\ : LocalMux
    port map (
            O => \N__4000\,
            I => \N__3997\
        );

    \I__763\ : Span12Mux_s9_v
    port map (
            O => \N__3997\,
            I => \N__3994\
        );

    \I__762\ : Span12Mux_h
    port map (
            O => \N__3994\,
            I => \N__3991\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__3991\,
            I => \un1_D_UU_040_7\
        );

    \I__760\ : InMux
    port map (
            O => \N__3988\,
            I => \N__3985\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__3982\,
            I => \N__3979\
        );

    \I__757\ : Sp12to4
    port map (
            O => \N__3979\,
            I => \N__3976\
        );

    \I__756\ : Span12Mux_h
    port map (
            O => \N__3976\,
            I => \N__3973\
        );

    \I__755\ : Odrv12
    port map (
            O => \N__3973\,
            I => \D_LL_AMIGA_in_3\
        );

    \I__754\ : IoInMux
    port map (
            O => \N__3970\,
            I => \N__3967\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3967\,
            I => \N__3964\
        );

    \I__752\ : IoSpan4Mux
    port map (
            O => \N__3964\,
            I => \N__3961\
        );

    \I__751\ : Sp12to4
    port map (
            O => \N__3961\,
            I => \N__3958\
        );

    \I__750\ : Span12Mux_s7_v
    port map (
            O => \N__3958\,
            I => \N__3955\
        );

    \I__749\ : Odrv12
    port map (
            O => \N__3955\,
            I => \un1_D_LL_AMIGA_3\
        );

    \I__748\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3949\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__3949\,
            I => \N__3946\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__3946\,
            I => \N__3943\
        );

    \I__745\ : Sp12to4
    port map (
            O => \N__3943\,
            I => \N__3940\
        );

    \I__744\ : Span12Mux_h
    port map (
            O => \N__3940\,
            I => \N__3937\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__3937\,
            I => \D_LL_AMIGA_in_1\
        );

    \I__742\ : IoInMux
    port map (
            O => \N__3934\,
            I => \N__3931\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3931\,
            I => \N__3928\
        );

    \I__740\ : Span12Mux_s3_h
    port map (
            O => \N__3928\,
            I => \N__3925\
        );

    \I__739\ : Span12Mux_h
    port map (
            O => \N__3925\,
            I => \N__3922\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__3922\,
            I => \un1_D_LL_AMIGA_1\
        );

    \I__737\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3916\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__3916\,
            I => \N__3912\
        );

    \I__735\ : IoInMux
    port map (
            O => \N__3915\,
            I => \N__3909\
        );

    \I__734\ : Span12Mux_h
    port map (
            O => \N__3912\,
            I => \N__3906\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3909\,
            I => \N__3903\
        );

    \I__732\ : Odrv12
    port map (
            O => \N__3906\,
            I => \A_AMIGA_c_1\
        );

    \I__731\ : Odrv12
    port map (
            O => \N__3903\,
            I => \A_AMIGA_c_1\
        );

    \I__730\ : IoInMux
    port map (
            O => \N__3898\,
            I => \N__3894\
        );

    \I__729\ : InMux
    port map (
            O => \N__3897\,
            I => \N__3891\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3894\,
            I => \N__3888\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__3891\,
            I => \N__3885\
        );

    \I__726\ : Span4Mux_s3_h
    port map (
            O => \N__3888\,
            I => \N__3882\
        );

    \I__725\ : Sp12to4
    port map (
            O => \N__3885\,
            I => \N__3879\
        );

    \I__724\ : Sp12to4
    port map (
            O => \N__3882\,
            I => \N__3876\
        );

    \I__723\ : Span12Mux_v
    port map (
            O => \N__3879\,
            I => \N__3873\
        );

    \I__722\ : Span12Mux_v
    port map (
            O => \N__3876\,
            I => \N__3870\
        );

    \I__721\ : Span12Mux_v
    port map (
            O => \N__3873\,
            I => \N__3865\
        );

    \I__720\ : Span12Mux_h
    port map (
            O => \N__3870\,
            I => \N__3865\
        );

    \I__719\ : Span12Mux_h
    port map (
            O => \N__3865\,
            I => \N__3862\
        );

    \I__718\ : Odrv12
    port map (
            O => \N__3862\,
            I => \D_LL_040_in_1\
        );

    \I__717\ : InMux
    port map (
            O => \N__3859\,
            I => \N__3856\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__3856\,
            I => \N__3853\
        );

    \I__715\ : Span4Mux_h
    port map (
            O => \N__3853\,
            I => \N__3850\
        );

    \I__714\ : Span4Mux_h
    port map (
            O => \N__3850\,
            I => \N__3847\
        );

    \I__713\ : Sp12to4
    port map (
            O => \N__3847\,
            I => \N__3844\
        );

    \I__712\ : Span12Mux_v
    port map (
            O => \N__3844\,
            I => \N__3841\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__3841\,
            I => \D_UM_040_in_1\
        );

    \I__710\ : IoInMux
    port map (
            O => \N__3838\,
            I => \N__3835\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__3835\,
            I => \N__3832\
        );

    \I__708\ : IoSpan4Mux
    port map (
            O => \N__3832\,
            I => \N__3829\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__3829\,
            I => \N__3826\
        );

    \I__706\ : Span12Mux_s6_h
    port map (
            O => \N__3826\,
            I => \N__3823\
        );

    \I__705\ : Odrv12
    port map (
            O => \N__3823\,
            I => \un1_D_UM_040_1\
        );

    \I__704\ : IoInMux
    port map (
            O => \N__3820\,
            I => \N__3817\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__3817\,
            I => \N__3814\
        );

    \I__702\ : IoSpan4Mux
    port map (
            O => \N__3814\,
            I => \N__3811\
        );

    \I__701\ : IoSpan4Mux
    port map (
            O => \N__3811\,
            I => \N__3808\
        );

    \I__700\ : Span4Mux_s2_v
    port map (
            O => \N__3808\,
            I => \N__3805\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__3805\,
            I => \N__3802\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__3802\,
            I => \LBENn_c_i\
        );

    \I__697\ : IoInMux
    port map (
            O => \N__3799\,
            I => \N__3796\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__3796\,
            I => \N__3793\
        );

    \I__695\ : Span4Mux_s3_h
    port map (
            O => \N__3793\,
            I => \N__3789\
        );

    \I__694\ : InMux
    port map (
            O => \N__3792\,
            I => \N__3786\
        );

    \I__693\ : Sp12to4
    port map (
            O => \N__3789\,
            I => \N__3783\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__3786\,
            I => \N__3780\
        );

    \I__691\ : Span12Mux_v
    port map (
            O => \N__3783\,
            I => \N__3777\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__3780\,
            I => \N__3774\
        );

    \I__689\ : Span12Mux_h
    port map (
            O => \N__3777\,
            I => \N__3769\
        );

    \I__688\ : Span12Mux_v
    port map (
            O => \N__3774\,
            I => \N__3769\
        );

    \I__687\ : Span12Mux_h
    port map (
            O => \N__3769\,
            I => \N__3766\
        );

    \I__686\ : Span12Mux_v
    port map (
            O => \N__3766\,
            I => \N__3763\
        );

    \I__685\ : Odrv12
    port map (
            O => \N__3763\,
            I => \D_LM_040_in_1\
        );

    \I__684\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3757\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__682\ : Sp12to4
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__681\ : Span12Mux_v
    port map (
            O => \N__3751\,
            I => \N__3748\
        );

    \I__680\ : Span12Mux_h
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__679\ : Odrv12
    port map (
            O => \N__3745\,
            I => \D_UU_040_in_1\
        );

    \I__678\ : IoInMux
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3739\,
            I => \N__3736\
        );

    \I__676\ : Span12Mux_s2_h
    port map (
            O => \N__3736\,
            I => \N__3733\
        );

    \I__675\ : Span12Mux_h
    port map (
            O => \N__3733\,
            I => \N__3730\
        );

    \I__674\ : Odrv12
    port map (
            O => \N__3730\,
            I => \un1_D_UU_040_1\
        );

    \I__673\ : IoInMux
    port map (
            O => \N__3727\,
            I => \N__3724\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__3724\,
            I => \N__3721\
        );

    \I__671\ : Span4Mux_s1_h
    port map (
            O => \N__3721\,
            I => \N__3718\
        );

    \I__670\ : Sp12to4
    port map (
            O => \N__3718\,
            I => \N__3714\
        );

    \I__669\ : InMux
    port map (
            O => \N__3717\,
            I => \N__3711\
        );

    \I__668\ : Span12Mux_v
    port map (
            O => \N__3714\,
            I => \N__3708\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__3711\,
            I => \N__3705\
        );

    \I__666\ : Span12Mux_h
    port map (
            O => \N__3708\,
            I => \N__3702\
        );

    \I__665\ : Span12Mux_h
    port map (
            O => \N__3705\,
            I => \N__3699\
        );

    \I__664\ : Span12Mux_h
    port map (
            O => \N__3702\,
            I => \N__3694\
        );

    \I__663\ : Span12Mux_v
    port map (
            O => \N__3699\,
            I => \N__3694\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__3694\,
            I => \D_LM_040_in_4\
        );

    \I__661\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__3688\,
            I => \N__3685\
        );

    \I__659\ : Span4Mux_v
    port map (
            O => \N__3685\,
            I => \N__3682\
        );

    \I__658\ : Sp12to4
    port map (
            O => \N__3682\,
            I => \N__3679\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__3679\,
            I => \N__3676\
        );

    \I__656\ : Odrv12
    port map (
            O => \N__3676\,
            I => \D_UU_040_in_4\
        );

    \I__655\ : IoInMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__3670\,
            I => \N__3667\
        );

    \I__653\ : IoSpan4Mux
    port map (
            O => \N__3667\,
            I => \N__3664\
        );

    \I__652\ : IoSpan4Mux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__651\ : Span4Mux_s3_v
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__650\ : Odrv4
    port map (
            O => \N__3658\,
            I => \un1_D_UU_040_4\
        );

    \I__649\ : InMux
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__3652\,
            I => \N__3649\
        );

    \I__647\ : Span12Mux_v
    port map (
            O => \N__3649\,
            I => \N__3646\
        );

    \I__646\ : Span12Mux_h
    port map (
            O => \N__3646\,
            I => \N__3643\
        );

    \I__645\ : Odrv12
    port map (
            O => \N__3643\,
            I => \D_UU_040_in_2\
        );

    \I__644\ : InMux
    port map (
            O => \N__3640\,
            I => \N__3637\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3637\,
            I => \N__3633\
        );

    \I__642\ : IoInMux
    port map (
            O => \N__3636\,
            I => \N__3630\
        );

    \I__641\ : Span4Mux_h
    port map (
            O => \N__3633\,
            I => \N__3627\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3630\,
            I => \N__3624\
        );

    \I__639\ : Span4Mux_h
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__638\ : Span12Mux_s9_h
    port map (
            O => \N__3624\,
            I => \N__3618\
        );

    \I__637\ : Sp12to4
    port map (
            O => \N__3621\,
            I => \N__3615\
        );

    \I__636\ : Span12Mux_h
    port map (
            O => \N__3618\,
            I => \N__3610\
        );

    \I__635\ : Span12Mux_v
    port map (
            O => \N__3615\,
            I => \N__3610\
        );

    \I__634\ : Span12Mux_v
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__633\ : Odrv12
    port map (
            O => \N__3607\,
            I => \D_LM_040_in_2\
        );

    \I__632\ : IoInMux
    port map (
            O => \N__3604\,
            I => \N__3601\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3601\,
            I => \N__3598\
        );

    \I__630\ : Span4Mux_s2_v
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__629\ : Span4Mux_v
    port map (
            O => \N__3595\,
            I => \N__3592\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__627\ : Odrv12
    port map (
            O => \N__3589\,
            I => \un1_D_UU_040_2\
        );

    \I__626\ : InMux
    port map (
            O => \N__3586\,
            I => \N__3583\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3583\,
            I => \N__3580\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__3580\,
            I => \N__3577\
        );

    \I__623\ : Sp12to4
    port map (
            O => \N__3577\,
            I => \N__3574\
        );

    \I__622\ : Span12Mux_h
    port map (
            O => \N__3574\,
            I => \N__3571\
        );

    \I__621\ : Odrv12
    port map (
            O => \N__3571\,
            I => \D_LL_AMIGA_in_2\
        );

    \I__620\ : IoInMux
    port map (
            O => \N__3568\,
            I => \N__3565\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3565\,
            I => \N__3562\
        );

    \I__618\ : Span12Mux_s4_h
    port map (
            O => \N__3562\,
            I => \N__3559\
        );

    \I__617\ : Span12Mux_h
    port map (
            O => \N__3559\,
            I => \N__3556\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__3556\,
            I => \un1_D_LL_AMIGA_2\
        );

    \I__615\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3550\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3550\,
            I => \N__3547\
        );

    \I__613\ : Span12Mux_v
    port map (
            O => \N__3547\,
            I => \N__3544\
        );

    \I__612\ : Span12Mux_h
    port map (
            O => \N__3544\,
            I => \N__3541\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__3541\,
            I => \D_LL_AMIGA_in_4\
        );

    \I__610\ : IoInMux
    port map (
            O => \N__3538\,
            I => \N__3535\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3535\,
            I => \N__3532\
        );

    \I__608\ : IoSpan4Mux
    port map (
            O => \N__3532\,
            I => \N__3529\
        );

    \I__607\ : Span4Mux_s2_h
    port map (
            O => \N__3529\,
            I => \N__3526\
        );

    \I__606\ : Sp12to4
    port map (
            O => \N__3526\,
            I => \N__3523\
        );

    \I__605\ : Span12Mux_h
    port map (
            O => \N__3523\,
            I => \N__3520\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__3520\,
            I => \un1_D_LL_AMIGA_4\
        );

    \I__603\ : InMux
    port map (
            O => \N__3517\,
            I => \N__3514\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3514\,
            I => \N__3511\
        );

    \I__601\ : Span12Mux_v
    port map (
            O => \N__3511\,
            I => \N__3508\
        );

    \I__600\ : Span12Mux_h
    port map (
            O => \N__3508\,
            I => \N__3505\
        );

    \I__599\ : Odrv12
    port map (
            O => \N__3505\,
            I => \D_LL_AMIGA_in_6\
        );

    \I__598\ : IoInMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__3499\,
            I => \N__3496\
        );

    \I__596\ : Span4Mux_s0_h
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__595\ : Span4Mux_h
    port map (
            O => \N__3493\,
            I => \N__3490\
        );

    \I__594\ : Sp12to4
    port map (
            O => \N__3490\,
            I => \N__3487\
        );

    \I__593\ : Span12Mux_s9_v
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__592\ : Span12Mux_h
    port map (
            O => \N__3484\,
            I => \N__3481\
        );

    \I__591\ : Odrv12
    port map (
            O => \N__3481\,
            I => \un1_D_LL_AMIGA_6\
        );

    \I__590\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3475\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__3472\,
            I => \N__3469\
        );

    \I__587\ : Sp12to4
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__586\ : Span12Mux_h
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__585\ : Odrv12
    port map (
            O => \N__3463\,
            I => \D_LM_AMIGA_in_0\
        );

    \I__584\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3457\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__3457\,
            I => \N__3454\
        );

    \I__582\ : Span4Mux_h
    port map (
            O => \N__3454\,
            I => \N__3451\
        );

    \I__581\ : Sp12to4
    port map (
            O => \N__3451\,
            I => \N__3448\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__3448\,
            I => \D_LM_AMIGA_in_2\
        );

    \I__579\ : IoInMux
    port map (
            O => \N__3445\,
            I => \N__3442\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3442\,
            I => \N__3439\
        );

    \I__577\ : Span12Mux_s6_h
    port map (
            O => \N__3439\,
            I => \N__3436\
        );

    \I__576\ : Span12Mux_v
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__3433\,
            I => \un1_D_LM_AMIGA_2\
        );

    \I__574\ : IoInMux
    port map (
            O => \N__3430\,
            I => \N__3427\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3427\,
            I => \N__3423\
        );

    \I__572\ : InMux
    port map (
            O => \N__3426\,
            I => \N__3420\
        );

    \I__571\ : IoSpan4Mux
    port map (
            O => \N__3423\,
            I => \N__3417\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3420\,
            I => \N__3414\
        );

    \I__569\ : Span4Mux_s3_h
    port map (
            O => \N__3417\,
            I => \N__3411\
        );

    \I__568\ : Span4Mux_h
    port map (
            O => \N__3414\,
            I => \N__3408\
        );

    \I__567\ : Sp12to4
    port map (
            O => \N__3411\,
            I => \N__3405\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__3408\,
            I => \N__3402\
        );

    \I__565\ : Span12Mux_v
    port map (
            O => \N__3405\,
            I => \N__3399\
        );

    \I__564\ : Span12Mux_v
    port map (
            O => \N__3402\,
            I => \N__3396\
        );

    \I__563\ : Span12Mux_h
    port map (
            O => \N__3399\,
            I => \N__3391\
        );

    \I__562\ : Span12Mux_v
    port map (
            O => \N__3396\,
            I => \N__3391\
        );

    \I__561\ : Span12Mux_h
    port map (
            O => \N__3391\,
            I => \N__3388\
        );

    \I__560\ : Odrv12
    port map (
            O => \N__3388\,
            I => \D_LL_040_in_7\
        );

    \I__559\ : InMux
    port map (
            O => \N__3385\,
            I => \N__3382\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__3382\,
            I => \N__3379\
        );

    \I__557\ : Span4Mux_v
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__556\ : Span4Mux_v
    port map (
            O => \N__3376\,
            I => \N__3373\
        );

    \I__555\ : Sp12to4
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__554\ : Span12Mux_h
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__553\ : Odrv12
    port map (
            O => \N__3367\,
            I => \D_UM_040_in_7\
        );

    \I__552\ : IoInMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3361\,
            I => \N__3358\
        );

    \I__550\ : IoSpan4Mux
    port map (
            O => \N__3358\,
            I => \N__3355\
        );

    \I__549\ : Span4Mux_s3_h
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__548\ : Span4Mux_h
    port map (
            O => \N__3352\,
            I => \N__3349\
        );

    \I__547\ : Span4Mux_h
    port map (
            O => \N__3349\,
            I => \N__3346\
        );

    \I__546\ : Odrv4
    port map (
            O => \N__3346\,
            I => \un1_D_UM_040_7\
        );

    \I__545\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3340\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3340\,
            I => \N__3337\
        );

    \I__543\ : Span4Mux_v
    port map (
            O => \N__3337\,
            I => \N__3334\
        );

    \I__542\ : Sp12to4
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__541\ : Span12Mux_h
    port map (
            O => \N__3331\,
            I => \N__3328\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3328\,
            I => \D_LL_AMIGA_in_0\
        );

    \I__539\ : IoInMux
    port map (
            O => \N__3325\,
            I => \N__3322\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__3322\,
            I => \N__3319\
        );

    \I__537\ : IoSpan4Mux
    port map (
            O => \N__3319\,
            I => \N__3316\
        );

    \I__536\ : IoSpan4Mux
    port map (
            O => \N__3316\,
            I => \N__3313\
        );

    \I__535\ : Span4Mux_s2_h
    port map (
            O => \N__3313\,
            I => \N__3310\
        );

    \I__534\ : Sp12to4
    port map (
            O => \N__3310\,
            I => \N__3307\
        );

    \I__533\ : Span12Mux_s9_h
    port map (
            O => \N__3307\,
            I => \N__3304\
        );

    \I__532\ : Odrv12
    port map (
            O => \N__3304\,
            I => \un1_D_LL_AMIGA_0\
        );

    \I__531\ : IoInMux
    port map (
            O => \N__3301\,
            I => \N__3298\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__3298\,
            I => \N__3295\
        );

    \I__529\ : Odrv12
    port map (
            O => \N__3295\,
            I => \LBENn_c_i_0\
        );

    \I__528\ : IoInMux
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3289\,
            I => \N__3286\
        );

    \I__526\ : Span12Mux_s6_v
    port map (
            O => \N__3286\,
            I => \N__3283\
        );

    \I__525\ : Odrv12
    port map (
            O => \N__3283\,
            I => \TSn_c\
        );

    \I__524\ : InMux
    port map (
            O => \N__3280\,
            I => \N__3277\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3277\,
            I => \N__3274\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__3274\,
            I => \N__3271\
        );

    \I__521\ : Sp12to4
    port map (
            O => \N__3271\,
            I => \N__3268\
        );

    \I__520\ : Span12Mux_h
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__519\ : Odrv12
    port map (
            O => \N__3265\,
            I => \D_LL_AMIGA_in_5\
        );

    \I__518\ : IoInMux
    port map (
            O => \N__3262\,
            I => \N__3259\
        );

    \I__517\ : LocalMux
    port map (
            O => \N__3259\,
            I => \N__3256\
        );

    \I__516\ : Span4Mux_s3_h
    port map (
            O => \N__3256\,
            I => \N__3253\
        );

    \I__515\ : Sp12to4
    port map (
            O => \N__3253\,
            I => \N__3250\
        );

    \I__514\ : Span12Mux_s11_v
    port map (
            O => \N__3250\,
            I => \N__3247\
        );

    \I__513\ : Span12Mux_h
    port map (
            O => \N__3247\,
            I => \N__3244\
        );

    \I__512\ : Odrv12
    port map (
            O => \N__3244\,
            I => \un1_D_LL_AMIGA_5\
        );

    \I__511\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3238\,
            I => \N__3235\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__3235\,
            I => \N__3232\
        );

    \I__508\ : Sp12to4
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__507\ : Span12Mux_h
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__506\ : Odrv12
    port map (
            O => \N__3226\,
            I => \D_LM_AMIGA_in_4\
        );

    \I__505\ : IoInMux
    port map (
            O => \N__3223\,
            I => \N__3220\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3220\,
            I => \N__3217\
        );

    \I__503\ : IoSpan4Mux
    port map (
            O => \N__3217\,
            I => \N__3214\
        );

    \I__502\ : IoSpan4Mux
    port map (
            O => \N__3214\,
            I => \N__3211\
        );

    \I__501\ : Span4Mux_s2_h
    port map (
            O => \N__3211\,
            I => \N__3208\
        );

    \I__500\ : Sp12to4
    port map (
            O => \N__3208\,
            I => \N__3205\
        );

    \I__499\ : Span12Mux_s11_h
    port map (
            O => \N__3205\,
            I => \N__3202\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__3202\,
            I => \un1_D_LM_AMIGA_4\
        );

    \I__497\ : InMux
    port map (
            O => \N__3199\,
            I => \N__3196\
        );

    \I__496\ : LocalMux
    port map (
            O => \N__3196\,
            I => \N__3193\
        );

    \I__495\ : Span12Mux_h
    port map (
            O => \N__3193\,
            I => \N__3190\
        );

    \I__494\ : Odrv12
    port map (
            O => \N__3190\,
            I => \D_UM_040_in_6\
        );

    \I__493\ : IoInMux
    port map (
            O => \N__3187\,
            I => \N__3184\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3184\,
            I => \N__3181\
        );

    \I__491\ : IoSpan4Mux
    port map (
            O => \N__3181\,
            I => \N__3177\
        );

    \I__490\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3174\
        );

    \I__489\ : IoSpan4Mux
    port map (
            O => \N__3177\,
            I => \N__3171\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3174\,
            I => \N__3168\
        );

    \I__487\ : Span4Mux_s2_h
    port map (
            O => \N__3171\,
            I => \N__3165\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__3168\,
            I => \N__3162\
        );

    \I__485\ : Sp12to4
    port map (
            O => \N__3165\,
            I => \N__3159\
        );

    \I__484\ : Sp12to4
    port map (
            O => \N__3162\,
            I => \N__3156\
        );

    \I__483\ : Span12Mux_h
    port map (
            O => \N__3159\,
            I => \N__3153\
        );

    \I__482\ : Span12Mux_h
    port map (
            O => \N__3156\,
            I => \N__3150\
        );

    \I__481\ : Span12Mux_h
    port map (
            O => \N__3153\,
            I => \N__3145\
        );

    \I__480\ : Span12Mux_v
    port map (
            O => \N__3150\,
            I => \N__3145\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__3145\,
            I => \D_LL_040_in_6\
        );

    \I__478\ : IoInMux
    port map (
            O => \N__3142\,
            I => \N__3139\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3139\,
            I => \N__3136\
        );

    \I__476\ : IoSpan4Mux
    port map (
            O => \N__3136\,
            I => \N__3133\
        );

    \I__475\ : Sp12to4
    port map (
            O => \N__3133\,
            I => \N__3130\
        );

    \I__474\ : Span12Mux_s6_h
    port map (
            O => \N__3130\,
            I => \N__3127\
        );

    \I__473\ : Span12Mux_v
    port map (
            O => \N__3127\,
            I => \N__3124\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__3124\,
            I => \un1_D_UM_040_6\
        );

    \I__471\ : IoInMux
    port map (
            O => \N__3121\,
            I => \N__3118\
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3118\,
            I => \N__3114\
        );

    \I__469\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3111\
        );

    \I__468\ : IoSpan4Mux
    port map (
            O => \N__3114\,
            I => \N__3108\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__3111\,
            I => \N__3105\
        );

    \I__466\ : Span4Mux_s2_h
    port map (
            O => \N__3108\,
            I => \N__3102\
        );

    \I__465\ : Span4Mux_v
    port map (
            O => \N__3105\,
            I => \N__3099\
        );

    \I__464\ : Sp12to4
    port map (
            O => \N__3102\,
            I => \N__3096\
        );

    \I__463\ : Sp12to4
    port map (
            O => \N__3099\,
            I => \N__3093\
        );

    \I__462\ : Span12Mux_h
    port map (
            O => \N__3096\,
            I => \N__3088\
        );

    \I__461\ : Span12Mux_v
    port map (
            O => \N__3093\,
            I => \N__3088\
        );

    \I__460\ : Span12Mux_h
    port map (
            O => \N__3088\,
            I => \N__3085\
        );

    \I__459\ : Odrv12
    port map (
            O => \N__3085\,
            I => \D_LL_040_in_2\
        );

    \I__458\ : InMux
    port map (
            O => \N__3082\,
            I => \N__3079\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3079\,
            I => \N__3076\
        );

    \I__456\ : Span12Mux_h
    port map (
            O => \N__3076\,
            I => \N__3073\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__3073\,
            I => \D_UM_040_in_2\
        );

    \I__454\ : IoInMux
    port map (
            O => \N__3070\,
            I => \N__3067\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__3067\,
            I => \N__3064\
        );

    \I__452\ : Span4Mux_s3_h
    port map (
            O => \N__3064\,
            I => \N__3061\
        );

    \I__451\ : Span4Mux_v
    port map (
            O => \N__3061\,
            I => \N__3058\
        );

    \I__450\ : Sp12to4
    port map (
            O => \N__3058\,
            I => \N__3055\
        );

    \I__449\ : Odrv12
    port map (
            O => \N__3055\,
            I => \un1_D_UM_040_2\
        );

    \I__448\ : InMux
    port map (
            O => \N__3052\,
            I => \N__3049\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3049\,
            I => \N__3046\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__3046\,
            I => \N__3043\
        );

    \I__445\ : Sp12to4
    port map (
            O => \N__3043\,
            I => \N__3040\
        );

    \I__444\ : Odrv12
    port map (
            O => \N__3040\,
            I => \D_LM_AMIGA_in_5\
        );

    \I__443\ : IoInMux
    port map (
            O => \N__3037\,
            I => \N__3034\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3034\,
            I => \N__3031\
        );

    \I__441\ : IoSpan4Mux
    port map (
            O => \N__3031\,
            I => \N__3028\
        );

    \I__440\ : Span4Mux_s2_h
    port map (
            O => \N__3028\,
            I => \N__3025\
        );

    \I__439\ : Span4Mux_v
    port map (
            O => \N__3025\,
            I => \N__3022\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__3022\,
            I => \N__3019\
        );

    \I__437\ : Span12Mux_s11_h
    port map (
            O => \N__3019\,
            I => \N__3016\
        );

    \I__436\ : Odrv12
    port map (
            O => \N__3016\,
            I => \un1_D_LM_AMIGA_5\
        );

    \I__435\ : InMux
    port map (
            O => \N__3013\,
            I => \N__3010\
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3010\,
            I => \N__3007\
        );

    \I__433\ : Span4Mux_h
    port map (
            O => \N__3007\,
            I => \N__3004\
        );

    \I__432\ : Span4Mux_v
    port map (
            O => \N__3004\,
            I => \N__3001\
        );

    \I__431\ : Sp12to4
    port map (
            O => \N__3001\,
            I => \N__2998\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__2998\,
            I => \D_LM_AMIGA_in_6\
        );

    \I__429\ : IoInMux
    port map (
            O => \N__2995\,
            I => \N__2992\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__2992\,
            I => \N__2989\
        );

    \I__427\ : Span12Mux_s2_h
    port map (
            O => \N__2989\,
            I => \N__2986\
        );

    \I__426\ : Span12Mux_h
    port map (
            O => \N__2986\,
            I => \N__2983\
        );

    \I__425\ : Odrv12
    port map (
            O => \N__2983\,
            I => \un1_D_LM_AMIGA_6\
        );

    \I__424\ : InMux
    port map (
            O => \N__2980\,
            I => \N__2976\
        );

    \I__423\ : IoInMux
    port map (
            O => \N__2979\,
            I => \N__2973\
        );

    \I__422\ : LocalMux
    port map (
            O => \N__2976\,
            I => \N__2970\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__2973\,
            I => \N__2967\
        );

    \I__420\ : Span4Mux_v
    port map (
            O => \N__2970\,
            I => \N__2964\
        );

    \I__419\ : Span4Mux_s2_h
    port map (
            O => \N__2967\,
            I => \N__2961\
        );

    \I__418\ : Sp12to4
    port map (
            O => \N__2964\,
            I => \N__2958\
        );

    \I__417\ : Span4Mux_v
    port map (
            O => \N__2961\,
            I => \N__2955\
        );

    \I__416\ : Span12Mux_h
    port map (
            O => \N__2958\,
            I => \N__2952\
        );

    \I__415\ : Sp12to4
    port map (
            O => \N__2955\,
            I => \N__2949\
        );

    \I__414\ : Span12Mux_v
    port map (
            O => \N__2952\,
            I => \N__2946\
        );

    \I__413\ : Span12Mux_s11_h
    port map (
            O => \N__2949\,
            I => \N__2943\
        );

    \I__412\ : Span12Mux_v
    port map (
            O => \N__2946\,
            I => \N__2938\
        );

    \I__411\ : Span12Mux_h
    port map (
            O => \N__2943\,
            I => \N__2938\
        );

    \I__410\ : Odrv12
    port map (
            O => \N__2938\,
            I => \D_LL_040_in_3\
        );

    \I__409\ : InMux
    port map (
            O => \N__2935\,
            I => \N__2932\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__2932\,
            I => \N__2929\
        );

    \I__407\ : Sp12to4
    port map (
            O => \N__2929\,
            I => \N__2926\
        );

    \I__406\ : Span12Mux_v
    port map (
            O => \N__2926\,
            I => \N__2923\
        );

    \I__405\ : Span12Mux_h
    port map (
            O => \N__2923\,
            I => \N__2920\
        );

    \I__404\ : Odrv12
    port map (
            O => \N__2920\,
            I => \D_UM_040_in_3\
        );

    \I__403\ : IoInMux
    port map (
            O => \N__2917\,
            I => \N__2914\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__2914\,
            I => \N__2911\
        );

    \I__401\ : IoSpan4Mux
    port map (
            O => \N__2911\,
            I => \N__2908\
        );

    \I__400\ : Span4Mux_s3_h
    port map (
            O => \N__2908\,
            I => \N__2905\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__2905\,
            I => \N__2902\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__2902\,
            I => \N__2899\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__2899\,
            I => \un1_D_UM_040_3\
        );

    \I__396\ : IoInMux
    port map (
            O => \N__2896\,
            I => \N__2893\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2893\,
            I => \N__2888\
        );

    \I__394\ : IoInMux
    port map (
            O => \N__2892\,
            I => \N__2883\
        );

    \I__393\ : IoInMux
    port map (
            O => \N__2891\,
            I => \N__2883\
        );

    \I__392\ : Span4Mux_s0_v
    port map (
            O => \N__2888\,
            I => \N__2879\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2883\,
            I => \N__2876\
        );

    \I__390\ : IoInMux
    port map (
            O => \N__2882\,
            I => \N__2873\
        );

    \I__389\ : Span4Mux_h
    port map (
            O => \N__2879\,
            I => \N__2870\
        );

    \I__388\ : Span4Mux_s0_v
    port map (
            O => \N__2876\,
            I => \N__2867\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__2873\,
            I => \N__2864\
        );

    \I__386\ : Span4Mux_h
    port map (
            O => \N__2870\,
            I => \N__2859\
        );

    \I__385\ : Span4Mux_h
    port map (
            O => \N__2867\,
            I => \N__2859\
        );

    \I__384\ : Span12Mux_s7_h
    port map (
            O => \N__2864\,
            I => \N__2856\
        );

    \I__383\ : Span4Mux_v
    port map (
            O => \N__2859\,
            I => \N__2853\
        );

    \I__382\ : Span12Mux_h
    port map (
            O => \N__2856\,
            I => \N__2850\
        );

    \I__381\ : Span4Mux_v
    port map (
            O => \N__2853\,
            I => \N__2847\
        );

    \I__380\ : Odrv12
    port map (
            O => \N__2850\,
            I => \CONSTANT_ONE_NET\
        );

    \I__379\ : Odrv4
    port map (
            O => \N__2847\,
            I => \CONSTANT_ONE_NET\
        );

    \I__378\ : InMux
    port map (
            O => \N__2842\,
            I => \N__2839\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2839\,
            I => \N__2836\
        );

    \I__376\ : Span4Mux_v
    port map (
            O => \N__2836\,
            I => \N__2833\
        );

    \I__375\ : Span4Mux_h
    port map (
            O => \N__2833\,
            I => \N__2830\
        );

    \I__374\ : Sp12to4
    port map (
            O => \N__2830\,
            I => \N__2827\
        );

    \I__373\ : Span12Mux_h
    port map (
            O => \N__2827\,
            I => \N__2824\
        );

    \I__372\ : Odrv12
    port map (
            O => \N__2824\,
            I => \D_UU_040_in_6\
        );

    \I__371\ : IoInMux
    port map (
            O => \N__2821\,
            I => \N__2818\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__2818\,
            I => \N__2815\
        );

    \I__369\ : Span4Mux_s2_h
    port map (
            O => \N__2815\,
            I => \N__2811\
        );

    \I__368\ : InMux
    port map (
            O => \N__2814\,
            I => \N__2808\
        );

    \I__367\ : Span4Mux_v
    port map (
            O => \N__2811\,
            I => \N__2805\
        );

    \I__366\ : LocalMux
    port map (
            O => \N__2808\,
            I => \N__2802\
        );

    \I__365\ : Sp12to4
    port map (
            O => \N__2805\,
            I => \N__2799\
        );

    \I__364\ : Sp12to4
    port map (
            O => \N__2802\,
            I => \N__2796\
        );

    \I__363\ : Span12Mux_h
    port map (
            O => \N__2799\,
            I => \N__2791\
        );

    \I__362\ : Span12Mux_s11_v
    port map (
            O => \N__2796\,
            I => \N__2791\
        );

    \I__361\ : Span12Mux_h
    port map (
            O => \N__2791\,
            I => \N__2788\
        );

    \I__360\ : Odrv12
    port map (
            O => \N__2788\,
            I => \D_LM_040_in_6\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__2785\,
            I => \N__2782\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__2782\,
            I => \N__2779\
        );

    \I__357\ : IoSpan4Mux
    port map (
            O => \N__2779\,
            I => \N__2776\
        );

    \I__356\ : Sp12to4
    port map (
            O => \N__2776\,
            I => \N__2773\
        );

    \I__355\ : Span12Mux_s6_v
    port map (
            O => \N__2773\,
            I => \N__2770\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__2770\,
            I => \un1_D_UU_040_6\
        );

    \I__353\ : InMux
    port map (
            O => \N__2767\,
            I => \N__2764\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__2764\,
            I => \N__2761\
        );

    \I__351\ : Span4Mux_v
    port map (
            O => \N__2761\,
            I => \N__2758\
        );

    \I__350\ : Span4Mux_h
    port map (
            O => \N__2758\,
            I => \N__2755\
        );

    \I__349\ : Sp12to4
    port map (
            O => \N__2755\,
            I => \N__2752\
        );

    \I__348\ : Span12Mux_h
    port map (
            O => \N__2752\,
            I => \N__2749\
        );

    \I__347\ : Odrv12
    port map (
            O => \N__2749\,
            I => \D_UU_040_in_0\
        );

    \I__346\ : IoInMux
    port map (
            O => \N__2746\,
            I => \N__2742\
        );

    \I__345\ : InMux
    port map (
            O => \N__2745\,
            I => \N__2739\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2742\,
            I => \N__2736\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__2739\,
            I => \N__2733\
        );

    \I__342\ : IoSpan4Mux
    port map (
            O => \N__2736\,
            I => \N__2730\
        );

    \I__341\ : Span4Mux_v
    port map (
            O => \N__2733\,
            I => \N__2727\
        );

    \I__340\ : IoSpan4Mux
    port map (
            O => \N__2730\,
            I => \N__2724\
        );

    \I__339\ : Sp12to4
    port map (
            O => \N__2727\,
            I => \N__2721\
        );

    \I__338\ : Span4Mux_s2_h
    port map (
            O => \N__2724\,
            I => \N__2718\
        );

    \I__337\ : Span12Mux_h
    port map (
            O => \N__2721\,
            I => \N__2715\
        );

    \I__336\ : Sp12to4
    port map (
            O => \N__2718\,
            I => \N__2712\
        );

    \I__335\ : Span12Mux_v
    port map (
            O => \N__2715\,
            I => \N__2709\
        );

    \I__334\ : Span12Mux_h
    port map (
            O => \N__2712\,
            I => \N__2706\
        );

    \I__333\ : Span12Mux_v
    port map (
            O => \N__2709\,
            I => \N__2701\
        );

    \I__332\ : Span12Mux_h
    port map (
            O => \N__2706\,
            I => \N__2701\
        );

    \I__331\ : Odrv12
    port map (
            O => \N__2701\,
            I => \D_LM_040_in_0\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__2698\,
            I => \N__2695\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__2695\,
            I => \N__2692\
        );

    \I__328\ : IoSpan4Mux
    port map (
            O => \N__2692\,
            I => \N__2689\
        );

    \I__327\ : IoSpan4Mux
    port map (
            O => \N__2689\,
            I => \N__2686\
        );

    \I__326\ : Span4Mux_s3_v
    port map (
            O => \N__2686\,
            I => \N__2683\
        );

    \I__325\ : Odrv4
    port map (
            O => \N__2683\,
            I => \un1_D_UU_040_0\
        );

    \I__324\ : InMux
    port map (
            O => \N__2680\,
            I => \N__2677\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2677\,
            I => \N__2674\
        );

    \I__322\ : Span12Mux_v
    port map (
            O => \N__2674\,
            I => \N__2671\
        );

    \I__321\ : Span12Mux_h
    port map (
            O => \N__2671\,
            I => \N__2668\
        );

    \I__320\ : Odrv12
    port map (
            O => \N__2668\,
            I => \D_LM_AMIGA_in_3\
        );

    \I__319\ : IoInMux
    port map (
            O => \N__2665\,
            I => \N__2662\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__2662\,
            I => \N__2659\
        );

    \I__317\ : Span4Mux_s0_h
    port map (
            O => \N__2659\,
            I => \N__2656\
        );

    \I__316\ : Sp12to4
    port map (
            O => \N__2656\,
            I => \N__2653\
        );

    \I__315\ : Span12Mux_v
    port map (
            O => \N__2653\,
            I => \N__2650\
        );

    \I__314\ : Span12Mux_h
    port map (
            O => \N__2650\,
            I => \N__2647\
        );

    \I__313\ : Odrv12
    port map (
            O => \N__2647\,
            I => \un1_D_LM_AMIGA_3\
        );

    \I__312\ : IoInMux
    port map (
            O => \N__2644\,
            I => \N__2641\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2641\,
            I => \N__2638\
        );

    \I__310\ : Span4Mux_s0_v
    port map (
            O => \N__2638\,
            I => \N__2635\
        );

    \I__309\ : Sp12to4
    port map (
            O => \N__2635\,
            I => \N__2632\
        );

    \I__308\ : Span12Mux_h
    port map (
            O => \N__2632\,
            I => \N__2629\
        );

    \I__307\ : Span12Mux_v
    port map (
            O => \N__2629\,
            I => \N__2626\
        );

    \I__306\ : Span12Mux_v
    port map (
            O => \N__2626\,
            I => \N__2623\
        );

    \I__305\ : Odrv12
    port map (
            O => \N__2623\,
            I => \TAn_in\
        );

    \I__304\ : InMux
    port map (
            O => \N__2620\,
            I => \N__2617\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__2617\,
            I => \N__2614\
        );

    \I__302\ : Span12Mux_h
    port map (
            O => \N__2614\,
            I => \N__2611\
        );

    \I__301\ : Odrv12
    port map (
            O => \N__2611\,
            I => \A_040_c_1\
        );

    \I__300\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2605\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2605\,
            I => \N__2602\
        );

    \I__298\ : Span4Mux_h
    port map (
            O => \N__2602\,
            I => \N__2599\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__2599\,
            I => \N__2596\
        );

    \I__296\ : Odrv4
    port map (
            O => \N__2596\,
            I => \A_040_c_0\
        );

    \I__295\ : IoInMux
    port map (
            O => \N__2593\,
            I => \N__2590\
        );

    \I__294\ : LocalMux
    port map (
            O => \N__2590\,
            I => \N__2587\
        );

    \I__293\ : Span4Mux_s2_v
    port map (
            O => \N__2587\,
            I => \N__2584\
        );

    \I__292\ : Span4Mux_v
    port map (
            O => \N__2584\,
            I => \N__2581\
        );

    \I__291\ : Odrv4
    port map (
            O => \N__2581\,
            I => \A_AMIGA_c_0\
        );

    \I__290\ : IoInMux
    port map (
            O => \N__2578\,
            I => \N__2575\
        );

    \I__289\ : LocalMux
    port map (
            O => \N__2575\,
            I => \N__2569\
        );

    \I__288\ : IoInMux
    port map (
            O => \N__2574\,
            I => \N__2566\
        );

    \I__287\ : IoInMux
    port map (
            O => \N__2573\,
            I => \N__2563\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2572\,
            I => \N__2560\
        );

    \I__285\ : IoSpan4Mux
    port map (
            O => \N__2569\,
            I => \N__2549\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__2566\,
            I => \N__2549\
        );

    \I__283\ : LocalMux
    port map (
            O => \N__2563\,
            I => \N__2549\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2560\,
            I => \N__2549\
        );

    \I__281\ : IoInMux
    port map (
            O => \N__2559\,
            I => \N__2546\
        );

    \I__280\ : IoInMux
    port map (
            O => \N__2558\,
            I => \N__2543\
        );

    \I__279\ : IoSpan4Mux
    port map (
            O => \N__2549\,
            I => \N__2535\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__2546\,
            I => \N__2535\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2543\,
            I => \N__2535\
        );

    \I__276\ : IoInMux
    port map (
            O => \N__2542\,
            I => \N__2532\
        );

    \I__275\ : IoSpan4Mux
    port map (
            O => \N__2535\,
            I => \N__2526\
        );

    \I__274\ : LocalMux
    port map (
            O => \N__2532\,
            I => \N__2523\
        );

    \I__273\ : IoInMux
    port map (
            O => \N__2531\,
            I => \N__2520\
        );

    \I__272\ : IoInMux
    port map (
            O => \N__2530\,
            I => \N__2517\
        );

    \I__271\ : IoInMux
    port map (
            O => \N__2529\,
            I => \N__2514\
        );

    \I__270\ : IoSpan4Mux
    port map (
            O => \N__2526\,
            I => \N__2496\
        );

    \I__269\ : IoSpan4Mux
    port map (
            O => \N__2523\,
            I => \N__2496\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2520\,
            I => \N__2496\
        );

    \I__267\ : LocalMux
    port map (
            O => \N__2517\,
            I => \N__2496\
        );

    \I__266\ : LocalMux
    port map (
            O => \N__2514\,
            I => \N__2496\
        );

    \I__265\ : IoInMux
    port map (
            O => \N__2513\,
            I => \N__2493\
        );

    \I__264\ : IoInMux
    port map (
            O => \N__2512\,
            I => \N__2490\
        );

    \I__263\ : IoInMux
    port map (
            O => \N__2511\,
            I => \N__2485\
        );

    \I__262\ : IoInMux
    port map (
            O => \N__2510\,
            I => \N__2482\
        );

    \I__261\ : IoInMux
    port map (
            O => \N__2509\,
            I => \N__2479\
        );

    \I__260\ : IoInMux
    port map (
            O => \N__2508\,
            I => \N__2476\
        );

    \I__259\ : IoInMux
    port map (
            O => \N__2507\,
            I => \N__2469\
        );

    \I__258\ : IoSpan4Mux
    port map (
            O => \N__2496\,
            I => \N__2460\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__2493\,
            I => \N__2460\
        );

    \I__256\ : LocalMux
    port map (
            O => \N__2490\,
            I => \N__2460\
        );

    \I__255\ : IoInMux
    port map (
            O => \N__2489\,
            I => \N__2457\
        );

    \I__254\ : IoInMux
    port map (
            O => \N__2488\,
            I => \N__2454\
        );

    \I__253\ : LocalMux
    port map (
            O => \N__2485\,
            I => \N__2440\
        );

    \I__252\ : LocalMux
    port map (
            O => \N__2482\,
            I => \N__2440\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2479\,
            I => \N__2440\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2476\,
            I => \N__2440\
        );

    \I__249\ : IoInMux
    port map (
            O => \N__2475\,
            I => \N__2437\
        );

    \I__248\ : IoInMux
    port map (
            O => \N__2474\,
            I => \N__2434\
        );

    \I__247\ : IoInMux
    port map (
            O => \N__2473\,
            I => \N__2431\
        );

    \I__246\ : IoInMux
    port map (
            O => \N__2472\,
            I => \N__2428\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__2469\,
            I => \N__2425\
        );

    \I__244\ : IoInMux
    port map (
            O => \N__2468\,
            I => \N__2422\
        );

    \I__243\ : IoInMux
    port map (
            O => \N__2467\,
            I => \N__2419\
        );

    \I__242\ : IoSpan4Mux
    port map (
            O => \N__2460\,
            I => \N__2412\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__2457\,
            I => \N__2412\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2454\,
            I => \N__2412\
        );

    \I__239\ : IoInMux
    port map (
            O => \N__2453\,
            I => \N__2409\
        );

    \I__238\ : IoInMux
    port map (
            O => \N__2452\,
            I => \N__2406\
        );

    \I__237\ : IoInMux
    port map (
            O => \N__2451\,
            I => \N__2403\
        );

    \I__236\ : IoInMux
    port map (
            O => \N__2450\,
            I => \N__2400\
        );

    \I__235\ : IoInMux
    port map (
            O => \N__2449\,
            I => \N__2397\
        );

    \I__234\ : IoSpan4Mux
    port map (
            O => \N__2440\,
            I => \N__2386\
        );

    \I__233\ : LocalMux
    port map (
            O => \N__2437\,
            I => \N__2386\
        );

    \I__232\ : LocalMux
    port map (
            O => \N__2434\,
            I => \N__2386\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__2431\,
            I => \N__2386\
        );

    \I__230\ : LocalMux
    port map (
            O => \N__2428\,
            I => \N__2371\
        );

    \I__229\ : IoSpan4Mux
    port map (
            O => \N__2425\,
            I => \N__2371\
        );

    \I__228\ : LocalMux
    port map (
            O => \N__2422\,
            I => \N__2371\
        );

    \I__227\ : LocalMux
    port map (
            O => \N__2419\,
            I => \N__2371\
        );

    \I__226\ : IoSpan4Mux
    port map (
            O => \N__2412\,
            I => \N__2371\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__2409\,
            I => \N__2371\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__2406\,
            I => \N__2371\
        );

    \I__223\ : LocalMux
    port map (
            O => \N__2403\,
            I => \N__2366\
        );

    \I__222\ : LocalMux
    port map (
            O => \N__2400\,
            I => \N__2366\
        );

    \I__221\ : LocalMux
    port map (
            O => \N__2397\,
            I => \N__2363\
        );

    \I__220\ : IoInMux
    port map (
            O => \N__2396\,
            I => \N__2360\
        );

    \I__219\ : IoInMux
    port map (
            O => \N__2395\,
            I => \N__2357\
        );

    \I__218\ : IoSpan4Mux
    port map (
            O => \N__2386\,
            I => \N__2354\
        );

    \I__217\ : IoSpan4Mux
    port map (
            O => \N__2371\,
            I => \N__2351\
        );

    \I__216\ : Span12Mux_s7_h
    port map (
            O => \N__2366\,
            I => \N__2348\
        );

    \I__215\ : Span12Mux_s9_h
    port map (
            O => \N__2363\,
            I => \N__2345\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__2360\,
            I => \N__2340\
        );

    \I__213\ : LocalMux
    port map (
            O => \N__2357\,
            I => \N__2340\
        );

    \I__212\ : Span4Mux_s1_v
    port map (
            O => \N__2354\,
            I => \N__2337\
        );

    \I__211\ : Span4Mux_s3_h
    port map (
            O => \N__2351\,
            I => \N__2334\
        );

    \I__210\ : Span12Mux_v
    port map (
            O => \N__2348\,
            I => \N__2331\
        );

    \I__209\ : Span12Mux_v
    port map (
            O => \N__2345\,
            I => \N__2326\
        );

    \I__208\ : Span12Mux_s9_h
    port map (
            O => \N__2340\,
            I => \N__2326\
        );

    \I__207\ : Span4Mux_v
    port map (
            O => \N__2337\,
            I => \N__2323\
        );

    \I__206\ : Span4Mux_h
    port map (
            O => \N__2334\,
            I => \N__2320\
        );

    \I__205\ : Odrv12
    port map (
            O => \N__2331\,
            I => \RnW_c_i\
        );

    \I__204\ : Odrv12
    port map (
            O => \N__2326\,
            I => \RnW_c_i\
        );

    \I__203\ : Odrv4
    port map (
            O => \N__2323\,
            I => \RnW_c_i\
        );

    \I__202\ : Odrv4
    port map (
            O => \N__2320\,
            I => \RnW_c_i\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            I => \N__4454\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            I => \N__4452\
        );

    \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            I => \N__4458\
        );

    \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            I => \N__4449\
        );

    \INVU111_CYCLE_SM.LW_CYCLEC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            I => \N__4451\
        );

    \INVU111_CYCLE_SM.CYCLE_STATE_1C\ : INV
    port map (
            O => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            I => \N__4453\
        );

    \INVU111_CYCLE_SM.TA_ENC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TA_ENC_net\,
            I => \N__4448\
        );

    \INVU111_CYCLE_SM.LW_CYCLE_STARTC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            I => \N__4450\
        );

    \INVU111_CYCLE_SM.TSnC\ : INV
    port map (
            O => \INVU111_CYCLE_SM.TSnC_net\,
            I => \N__5673\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNIK8GP_LC_3_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4396\,
            in1 => \N__2620\,
            in2 => \_gnd_net_\,
            in3 => \N__7272\,
            lcout => \A_AMIGA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIN15M_LC_3_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__2608\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7273\,
            lcout => \A_AMIGA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RnW_c_sbtinv_LC_6_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6041\,
            lcout => \RnW_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOROB2_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3117\,
            in1 => \N__4759\,
            in2 => \_gnd_net_\,
            in3 => \N__3082\,
            lcout => \un1_D_UM_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITNJF2_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3052\,
            in1 => \N__4859\,
            in2 => \_gnd_net_\,
            in3 => \N__6825\,
            lcout => \un1_D_LM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVPJF2_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4860\,
            in1 => \N__6554\,
            in2 => \_gnd_net_\,
            in3 => \N__3013\,
            lcout => \un1_D_LM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIQTOB2_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__2980\,
            in1 => \N__4869\,
            in2 => \_gnd_net_\,
            in3 => \N__2935\,
            lcout => \un1_D_UM_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI9PQV1_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4879\,
            in1 => \N__2842\,
            in2 => \_gnd_net_\,
            in3 => \N__2814\,
            lcout => \un1_D_UU_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNITCQV1_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2767\,
            in1 => \N__4880\,
            in2 => \_gnd_net_\,
            in3 => \N__2745\,
            lcout => \un1_D_UU_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIPJJF2_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__4830\,
            in2 => \_gnd_net_\,
            in3 => \N__2680\,
            lcout => \un1_D_LM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNINHJF2_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4829\,
            in1 => \N__5548\,
            in2 => \_gnd_net_\,
            in3 => \N__3460\,
            lcout => \un1_D_LM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI26PB2_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3426\,
            in1 => \N__4878\,
            in2 => \_gnd_net_\,
            in3 => \N__3385\,
            lcout => \un1_D_UM_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIA6UI2_LC_11_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3343\,
            in1 => \N__4855\,
            in2 => \_gnd_net_\,
            in3 => \N__6466\,
            lcout => \un1_D_LL_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \LBENn_c_sbtinv_LC_11_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5831\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \LBENn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TSn_LC_11_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__6094\,
            in1 => \_gnd_net_\,
            in2 => \N__5849\,
            in3 => \N__5146\,
            lcout => \TSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TSnC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKGUI2_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6772\,
            in1 => \N__4814\,
            in2 => \_gnd_net_\,
            in3 => \N__3280\,
            lcout => \un1_D_LL_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIRLJF2_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4818\,
            in1 => \N__6634\,
            in2 => \_gnd_net_\,
            in3 => \N__3241\,
            lcout => \un1_D_LM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI04PB2_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4817\,
            in1 => \N__3199\,
            in2 => \_gnd_net_\,
            in3 => \N__3180\,
            lcout => \un1_D_UM_040_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMPOB2_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3897\,
            in1 => \N__4870\,
            in2 => \_gnd_net_\,
            in3 => \N__3859\,
            lcout => \un1_D_UM_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \BUFENn_obuf_RNO_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5867\,
            lcout => \LBENn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIVEQV1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3792\,
            in1 => \N__4871\,
            in2 => \_gnd_net_\,
            in3 => \N__3760\,
            lcout => \un1_D_UU_040_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI5LQV1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3717\,
            in1 => \N__4882\,
            in2 => \_gnd_net_\,
            in3 => \N__3691\,
            lcout => \un1_D_UU_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1HQV1_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3655\,
            in1 => \N__4881\,
            in2 => \_gnd_net_\,
            in3 => \N__3640\,
            lcout => \un1_D_UU_040_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIEAUI2_LC_12_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6367\,
            in1 => \N__4815\,
            in2 => \_gnd_net_\,
            in3 => \N__3586\,
            lcout => \un1_D_LL_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIIEUI2_LC_12_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4816\,
            in1 => \N__7324\,
            in2 => \_gnd_net_\,
            in3 => \N__3553\,
            lcout => \un1_D_LL_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIMIUI2_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6415\,
            in1 => \N__4819\,
            in2 => \_gnd_net_\,
            in3 => \N__3517\,
            lcout => \un1_D_LL_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIJDJF2_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4760\,
            in1 => \N__6910\,
            in2 => \_gnd_net_\,
            in3 => \N__3478\,
            lcout => \un1_D_LM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIOKUI2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__6974\,
            in1 => \N__4761\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \un1_D_LL_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIKNOB2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4708\,
            in1 => \N__4311\,
            in2 => \_gnd_net_\,
            in3 => \N__4270\,
            lcout => \un1_D_UM_040_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNISVOB2_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__4856\,
            in1 => \N__4237\,
            in2 => \_gnd_net_\,
            in3 => \N__4216\,
            lcout => \un1_D_UM_040_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI7NQV1_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4146\,
            in1 => \N__4857\,
            in2 => \_gnd_net_\,
            in3 => \N__4105\,
            lcout => \un1_D_UU_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIBRQV1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4858\,
            in1 => \N__4056\,
            in2 => \_gnd_net_\,
            in3 => \N__4021\,
            lcout => \un1_D_UU_040_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIGCUI2_LC_13_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3988\,
            in1 => \N__4808\,
            in2 => \_gnd_net_\,
            in3 => \N__7123\,
            lcout => \un1_D_LL_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIC8UI2_LC_13_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5770\,
            in1 => \N__4807\,
            in2 => \_gnd_net_\,
            in3 => \N__3952\,
            lcout => \un1_D_LL_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIM3VM1_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__7263\,
            in1 => \N__5038\,
            in2 => \_gnd_net_\,
            in3 => \N__3919\,
            lcout => \U111_CYCLE_SM.FLIP\,
            ltout => \U111_CYCLE_SM.FLIP_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNILFJF2_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__4558\,
            in1 => \_gnd_net_\,
            in2 => \N__4546\,
            in3 => \N__5977\,
            lcout => \un1_D_LM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_THRU_LUT4_0_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5689\,
            lcout => \GB_BUFFER_CLK40_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK80_THRU_LUT4_0_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_CLK80_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011000000"
        )
    port map (
            in0 => \N__7189\,
            in1 => \N__5122\,
            in2 => \N__6148\,
            in3 => \N__5180\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_RNO_0_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101110"
        )
    port map (
            in0 => \N__6198\,
            in1 => \N__4386\,
            in2 => \N__5182\,
            in3 => \N__6247\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.A_OUT_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.A_OUT_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4399\,
            in3 => \N__6129\,
            lcout => \U111_CYCLE_SM.A_OUTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110011001"
        )
    port map (
            in0 => \N__6197\,
            in1 => \N__6246\,
            in2 => \_gnd_net_\,
            in3 => \N__5687\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_75_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__5139\,
            in1 => \N__6130\,
            in2 => \N__4375\,
            in3 => \N__4564\,
            lcout => \U111_CYCLE_SM.TS_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNO_0_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__6137\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_START_RNO_0_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5064\,
            in1 => \N__5037\,
            in2 => \N__5871\,
            in3 => \N__5138\,
            lcout => \U111_CYCLE_SM.un3_LW_CYCLE_START\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000011011100"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__6201\,
            in2 => \N__5903\,
            in3 => \N__6248\,
            lcout => \U111_CYCLE_SM.TA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.TA_ENC_net\,
            ce => 'H',
            sr => \N__5116\
        );

    \U111_CYCLE_SM.LW_TRANS_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__5104\,
            in1 => \N__5086\,
            in2 => \_gnd_net_\,
            in3 => \N__5068\,
            lcout => \U111_CYCLE_SM.LW_TRANS_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI1SJF2_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5625\,
            in1 => \N__4820\,
            in2 => \_gnd_net_\,
            in3 => \N__5020\,
            lcout => \un1_D_LM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNIU1PB2_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__4813\,
            in2 => \_gnd_net_\,
            in3 => \N__4933\,
            lcout => \un1_D_UM_040_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNI3JQV1_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4900\,
            in1 => \N__4812\,
            in2 => \_gnd_net_\,
            in3 => \N__4650\,
            lcout => \un1_D_UU_040_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNI4SHG_LC_14_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__5911\,
            in1 => \N__6275\,
            in2 => \_gnd_net_\,
            in3 => \N__5850\,
            lcout => \U111_CYCLE_SM_TBI_CPUn_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_1_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__6192\,
            in1 => \N__5479\,
            in2 => \N__6250\,
            in3 => \N__5647\,
            lcout => \U111_CYCLE_SM.TS_EN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CPU_READ_EN_i_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5478\,
            in1 => \N__6045\,
            in2 => \_gnd_net_\,
            in3 => \N__5866\,
            lcout => \CPU_READ_EN_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_1_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001000010100000"
        )
    port map (
            in0 => \N__6193\,
            in1 => \N__6282\,
            in2 => \N__6154\,
            in3 => \N__6249\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.CYCLE_STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_0_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5175\,
            in2 => \_gnd_net_\,
            in3 => \N__6241\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.A_OUT_0_sqmuxa_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010101000"
        )
    port map (
            in0 => \N__6152\,
            in1 => \N__5152\,
            in2 => \N__5185\,
            in3 => \N__6200\,
            lcout => \U111_CYCLE_SM.LW_CYCLEZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNO_0_0_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__6199\,
            in1 => \N__5176\,
            in2 => \_gnd_net_\,
            in3 => \N__5688\,
            lcout => OPEN,
            ltout => \U111_CYCLE_SM.N_97_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__6242\,
            in1 => \N__6301\,
            in2 => \N__5155\,
            in3 => \N__6147\,
            lcout => \U111_CYCLE_SM.CYCLE_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.LW_CYCLEC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.LW_CYCLE_RNO_1_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001001100"
        )
    port map (
            in0 => \N__6240\,
            in1 => \N__7188\,
            in2 => \N__6202\,
            in3 => \N__6302\,
            lcout => \U111_CYCLE_SM.LW_CYCLE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_2_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5547\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7045\,
            sr => \N__7005\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_7_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5621\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7045\,
            sr => \N__7005\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_1_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5973\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7045\,
            sr => \N__7005\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_1_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__5766\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UU_LATCHED_nesr_2C_net\,
            ce => \N__7045\,
            sr => \N__7005\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI0IN51_1_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7228\,
            in1 => \N__5983\,
            in2 => \_gnd_net_\,
            in3 => \N__5972\,
            lcout => \un1_D_UU_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TA_EN_RNIVCEG_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5904\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5878\,
            lcout => \TAn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIGP7L_1_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5753\,
            in1 => \N__5725\,
            in2 => \_gnd_net_\,
            in3 => \N__7227\,
            lcout => \un1_D_UM_AMIGA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.TS_EN_RNO_2_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5701\,
            in2 => \_gnd_net_\,
            in3 => \N__5686\,
            lcout => \U111_CYCLE_SM.TS_EN_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNICUN51_7_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7230\,
            in1 => \N__5635\,
            in2 => \_gnd_net_\,
            in3 => \N__5626\,
            lcout => \un1_D_UU_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI2KN51_2_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__5543\,
            in2 => \_gnd_net_\,
            in3 => \N__7229\,
            lcout => \un1_D_UU_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIEN7L_0_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6424\,
            in1 => \N__6459\,
            in2 => \_gnd_net_\,
            in3 => \N__7249\,
            lcout => \un1_D_UM_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIIR7L_2_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7250\,
            in1 => \N__6325\,
            in2 => \_gnd_net_\,
            in3 => \N__6360\,
            lcout => \un1_D_UM_AMIGA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIQ38L_6_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6373\,
            in1 => \N__6401\,
            in2 => \_gnd_net_\,
            in3 => \N__7248\,
            lcout => \un1_D_UM_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_0_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6458\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            ce => \N__7036\,
            sr => \N__7003\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_6_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6411\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            ce => \N__7036\,
            sr => \N__7003\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6359\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_0C_net\,
            ce => \N__7036\,
            sr => \N__7003\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIULFD_0_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6303\,
            in1 => \N__6239\,
            in2 => \_gnd_net_\,
            in3 => \N__6191\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1_0_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6153\,
            in2 => \N__6055\,
            in3 => \N__6037\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0\,
            ltout => \U111_CYCLE_SM.CYCLE_STATE_RNIGD9C1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.CYCLE_STATE_RNIE3PP1_0_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5992\,
            in3 => \N__5989\,
            lcout => \U111_CYCLE_SM.CYCLE_STATE_0_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_3_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7119\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7044\,
            sr => \N__7004\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_5_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6764\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7044\,
            sr => \N__7004\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_3_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6694\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7044\,
            sr => \N__7004\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_4_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6630\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7044\,
            sr => \N__7004\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_6_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6562\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_3C_net\,
            ce => \N__7044\,
            sr => \N__7004\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIO18L_5_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7231\,
            in1 => \N__6778\,
            in2 => \_gnd_net_\,
            in3 => \N__6771\,
            lcout => \un1_D_UM_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI4MN51_3_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7232\,
            in1 => \N__6700\,
            in2 => \_gnd_net_\,
            in3 => \N__6693\,
            lcout => \un1_D_UU_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI6ON51_4_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7233\,
            in1 => \N__6640\,
            in2 => \_gnd_net_\,
            in3 => \N__6629\,
            lcout => \un1_D_UU_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIASN51_6_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7262\,
            in1 => \N__6571\,
            in2 => \_gnd_net_\,
            in3 => \N__6561\,
            lcout => \un1_D_UU_AMIGA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIKT7L_3_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7112\,
            in1 => \N__7075\,
            in2 => \_gnd_net_\,
            in3 => \N__7261\,
            lcout => \un1_D_UM_AMIGA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_4_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7320\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__7043\,
            sr => \N__7006\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_5_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6841\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__7043\,
            sr => \N__7006\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_0_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6906\,
            lcout => \U111_CYCLE_SM.UU_LATCHEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__7043\,
            sr => \N__7006\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_7_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6976\,
            lcout => \U111_CYCLE_SM.UM_LATCHEDZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU111_CYCLE_SM.UM_LATCHED_nesr_4C_net\,
            ce => \N__7043\,
            sr => \N__7006\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIS58L_7_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7258\,
            in1 => \N__6982\,
            in2 => \_gnd_net_\,
            in3 => \N__6975\,
            lcout => \un1_D_UM_AMIGA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNIUFN51_0_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7260\,
            in1 => \N__6916\,
            in2 => \_gnd_net_\,
            in3 => \N__6905\,
            lcout => \un1_D_UU_AMIGA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UU_LATCHED_nesr_RNI8QN51_5_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6847\,
            in1 => \N__6837\,
            in2 => \_gnd_net_\,
            in3 => \N__7259\,
            lcout => \un1_D_UU_AMIGA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U111_CYCLE_SM.UM_LATCHED_nesr_RNIMV7L_4_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7330\,
            in1 => \N__7319\,
            in2 => \_gnd_net_\,
            in3 => \N__7257\,
            lcout => \un1_D_UM_AMIGA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

module U109_PCI_STATE_MACHINE (

    output PCICYCLEn, ADLATCH, ALATCH, PCIDIR

);

//DISABLE THE ADDRESS BUFFERS FOR NOW.

//ADDRESS DATA IS PASSED THROUGH LIVE DURING THE ADDRESS PHASE OF CPU DRIVEN CYCLES.
//FOR PCI DRIVEN DMA CYCLES, THE ADDRESS IS LATCHED DURING THE ADDRESS PHASE AND
//DRIVEN ON THE ADDRESS BUS OF THE AMIGAPCI.

assign PCICYCLEn = 1;
assign ADLATCH = 0;
assign ALATCH = 0; //WE DON'T ACTUALLY NEED THIS, BUT ITS THERE.
assign PCIDIR = 0;


endmodule

// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 13 2025 19:08:48

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "U712_TOP" view "INTERFACE"

module U712_TOP (
    SIZ,
    CMA,
    DRA,
    DA,
    A,
    DBRn,
    TSn,
    LMBEn,
    DMA_LATCH_EN,
    CLMBEn,
    AWEn,
    RESETn,
    CLK_EN,
    CASn,
    BANK0,
    CLK40B_OUT,
    VBENn,
    CUMBEn,
    CLKRAM,
    CLK40D_OUT,
    C3,
    ASn,
    UUBEn,
    LDSn,
    LATCH_CLK,
    CASUn,
    RAS1n,
    DRDDIR,
    DBDIR,
    UDSn,
    RnW,
    DRDENn,
    DBENn,
    BANK1,
    UMBEn,
    RAS0n,
    CUUBEn,
    CRCSn,
    CLLBEn,
    CLK40C_OUT,
    CASLn,
    TCIn,
    TBIn,
    RAMSPACEn,
    WEn,
    REGENn,
    LLBEn,
    CLK40_IN,
    REGSPACEn,
    RASn,
    AGNUS_REV,
    TACKn,
    C1);

    input [1:0] SIZ;
    output [10:0] CMA;
    input [9:0] DRA;
    output [2:0] DA;
    input [20:0] A;
    input DBRn;
    input TSn;
    output LMBEn;
    output DMA_LATCH_EN;
    output CLMBEn;
    input AWEn;
    input RESETn;
    output CLK_EN;
    output CASn;
    output BANK0;
    output CLK40B_OUT;
    output VBENn;
    output CUMBEn;
    output CLKRAM;
    output CLK40D_OUT;
    input C3;
    output ASn;
    output UUBEn;
    output LDSn;
    output LATCH_CLK;
    input CASUn;
    input RAS1n;
    output DRDDIR;
    output DBDIR;
    output UDSn;
    input RnW;
    output DRDENn;
    output DBENn;
    output BANK1;
    output UMBEn;
    input RAS0n;
    output CUUBEn;
    output CRCSn;
    output CLLBEn;
    output CLK40C_OUT;
    input CASLn;
    output TCIn;
    output TBIn;
    input RAMSPACEn;
    output WEn;
    output REGENn;
    output LLBEn;
    input CLK40_IN;
    input REGSPACEn;
    output RASn;
    input AGNUS_REV;
    output TACKn;
    input C1;

    wire N__12615;
    wire N__12614;
    wire N__12613;
    wire N__12606;
    wire N__12605;
    wire N__12604;
    wire N__12597;
    wire N__12596;
    wire N__12595;
    wire N__12588;
    wire N__12587;
    wire N__12586;
    wire N__12579;
    wire N__12578;
    wire N__12577;
    wire N__12570;
    wire N__12569;
    wire N__12568;
    wire N__12561;
    wire N__12560;
    wire N__12559;
    wire N__12552;
    wire N__12551;
    wire N__12550;
    wire N__12543;
    wire N__12542;
    wire N__12541;
    wire N__12534;
    wire N__12533;
    wire N__12532;
    wire N__12525;
    wire N__12524;
    wire N__12523;
    wire N__12516;
    wire N__12515;
    wire N__12514;
    wire N__12507;
    wire N__12506;
    wire N__12505;
    wire N__12498;
    wire N__12497;
    wire N__12496;
    wire N__12489;
    wire N__12488;
    wire N__12487;
    wire N__12480;
    wire N__12479;
    wire N__12478;
    wire N__12471;
    wire N__12470;
    wire N__12469;
    wire N__12462;
    wire N__12461;
    wire N__12460;
    wire N__12453;
    wire N__12452;
    wire N__12451;
    wire N__12444;
    wire N__12443;
    wire N__12442;
    wire N__12435;
    wire N__12434;
    wire N__12433;
    wire N__12426;
    wire N__12425;
    wire N__12424;
    wire N__12417;
    wire N__12416;
    wire N__12415;
    wire N__12408;
    wire N__12407;
    wire N__12406;
    wire N__12399;
    wire N__12398;
    wire N__12397;
    wire N__12390;
    wire N__12389;
    wire N__12388;
    wire N__12381;
    wire N__12380;
    wire N__12379;
    wire N__12372;
    wire N__12371;
    wire N__12370;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12354;
    wire N__12353;
    wire N__12352;
    wire N__12345;
    wire N__12344;
    wire N__12343;
    wire N__12336;
    wire N__12335;
    wire N__12334;
    wire N__12327;
    wire N__12326;
    wire N__12325;
    wire N__12318;
    wire N__12317;
    wire N__12316;
    wire N__12309;
    wire N__12308;
    wire N__12307;
    wire N__12300;
    wire N__12299;
    wire N__12298;
    wire N__12291;
    wire N__12290;
    wire N__12289;
    wire N__12282;
    wire N__12281;
    wire N__12280;
    wire N__12273;
    wire N__12272;
    wire N__12271;
    wire N__12264;
    wire N__12263;
    wire N__12262;
    wire N__12255;
    wire N__12254;
    wire N__12253;
    wire N__12246;
    wire N__12245;
    wire N__12244;
    wire N__12237;
    wire N__12236;
    wire N__12235;
    wire N__12228;
    wire N__12227;
    wire N__12226;
    wire N__12219;
    wire N__12218;
    wire N__12217;
    wire N__12210;
    wire N__12209;
    wire N__12208;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12192;
    wire N__12191;
    wire N__12190;
    wire N__12183;
    wire N__12182;
    wire N__12181;
    wire N__12174;
    wire N__12173;
    wire N__12172;
    wire N__12165;
    wire N__12164;
    wire N__12163;
    wire N__12156;
    wire N__12155;
    wire N__12154;
    wire N__12147;
    wire N__12146;
    wire N__12145;
    wire N__12138;
    wire N__12137;
    wire N__12136;
    wire N__12129;
    wire N__12128;
    wire N__12127;
    wire N__12120;
    wire N__12119;
    wire N__12118;
    wire N__12111;
    wire N__12110;
    wire N__12109;
    wire N__12102;
    wire N__12101;
    wire N__12100;
    wire N__12093;
    wire N__12092;
    wire N__12091;
    wire N__12084;
    wire N__12083;
    wire N__12082;
    wire N__12075;
    wire N__12074;
    wire N__12073;
    wire N__12066;
    wire N__12065;
    wire N__12064;
    wire N__12057;
    wire N__12056;
    wire N__12055;
    wire N__12048;
    wire N__12047;
    wire N__12046;
    wire N__12039;
    wire N__12038;
    wire N__12037;
    wire N__12030;
    wire N__12029;
    wire N__12028;
    wire N__12021;
    wire N__12020;
    wire N__12019;
    wire N__12012;
    wire N__12011;
    wire N__12010;
    wire N__12003;
    wire N__12002;
    wire N__12001;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11985;
    wire N__11984;
    wire N__11983;
    wire N__11976;
    wire N__11975;
    wire N__11974;
    wire N__11967;
    wire N__11966;
    wire N__11965;
    wire N__11958;
    wire N__11957;
    wire N__11956;
    wire N__11949;
    wire N__11948;
    wire N__11947;
    wire N__11940;
    wire N__11939;
    wire N__11938;
    wire N__11931;
    wire N__11930;
    wire N__11929;
    wire N__11922;
    wire N__11921;
    wire N__11920;
    wire N__11913;
    wire N__11912;
    wire N__11911;
    wire N__11904;
    wire N__11903;
    wire N__11902;
    wire N__11895;
    wire N__11894;
    wire N__11893;
    wire N__11886;
    wire N__11885;
    wire N__11884;
    wire N__11877;
    wire N__11876;
    wire N__11875;
    wire N__11868;
    wire N__11867;
    wire N__11866;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11850;
    wire N__11849;
    wire N__11848;
    wire N__11841;
    wire N__11840;
    wire N__11839;
    wire N__11832;
    wire N__11831;
    wire N__11830;
    wire N__11823;
    wire N__11822;
    wire N__11821;
    wire N__11814;
    wire N__11813;
    wire N__11812;
    wire N__11805;
    wire N__11804;
    wire N__11803;
    wire N__11796;
    wire N__11795;
    wire N__11794;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11778;
    wire N__11777;
    wire N__11776;
    wire N__11769;
    wire N__11768;
    wire N__11767;
    wire N__11750;
    wire N__11749;
    wire N__11748;
    wire N__11745;
    wire N__11744;
    wire N__11743;
    wire N__11738;
    wire N__11735;
    wire N__11732;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11707;
    wire N__11700;
    wire N__11697;
    wire N__11692;
    wire N__11687;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11677;
    wire N__11674;
    wire N__11671;
    wire N__11670;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11620;
    wire N__11615;
    wire N__11614;
    wire N__11613;
    wire N__11612;
    wire N__11611;
    wire N__11610;
    wire N__11609;
    wire N__11606;
    wire N__11599;
    wire N__11596;
    wire N__11591;
    wire N__11588;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11552;
    wire N__11551;
    wire N__11550;
    wire N__11549;
    wire N__11548;
    wire N__11547;
    wire N__11540;
    wire N__11535;
    wire N__11534;
    wire N__11531;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11510;
    wire N__11507;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11495;
    wire N__11492;
    wire N__11487;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11471;
    wire N__11470;
    wire N__11467;
    wire N__11466;
    wire N__11465;
    wire N__11464;
    wire N__11463;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11440;
    wire N__11437;
    wire N__11432;
    wire N__11429;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11411;
    wire N__11406;
    wire N__11403;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11380;
    wire N__11379;
    wire N__11376;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11362;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11350;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11337;
    wire N__11336;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11301;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11218;
    wire N__11217;
    wire N__11214;
    wire N__11211;
    wire N__11208;
    wire N__11207;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11195;
    wire N__11192;
    wire N__11187;
    wire N__11184;
    wire N__11179;
    wire N__11174;
    wire N__11173;
    wire N__11172;
    wire N__11169;
    wire N__11168;
    wire N__11165;
    wire N__11164;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11131;
    wire N__11126;
    wire N__11123;
    wire N__11118;
    wire N__11113;
    wire N__11110;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11089;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11046;
    wire N__11043;
    wire N__11038;
    wire N__11033;
    wire N__11030;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10999;
    wire N__10998;
    wire N__10997;
    wire N__10996;
    wire N__10995;
    wire N__10994;
    wire N__10991;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10983;
    wire N__10982;
    wire N__10981;
    wire N__10980;
    wire N__10979;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10954;
    wire N__10949;
    wire N__10946;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10938;
    wire N__10937;
    wire N__10936;
    wire N__10935;
    wire N__10934;
    wire N__10933;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10905;
    wire N__10902;
    wire N__10899;
    wire N__10896;
    wire N__10889;
    wire N__10886;
    wire N__10879;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10855;
    wire N__10852;
    wire N__10847;
    wire N__10846;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10832;
    wire N__10829;
    wire N__10824;
    wire N__10821;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10789;
    wire N__10788;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10768;
    wire N__10767;
    wire N__10766;
    wire N__10765;
    wire N__10764;
    wire N__10763;
    wire N__10762;
    wire N__10761;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10735;
    wire N__10734;
    wire N__10733;
    wire N__10732;
    wire N__10731;
    wire N__10730;
    wire N__10729;
    wire N__10726;
    wire N__10719;
    wire N__10716;
    wire N__10711;
    wire N__10708;
    wire N__10707;
    wire N__10704;
    wire N__10703;
    wire N__10702;
    wire N__10701;
    wire N__10700;
    wire N__10699;
    wire N__10698;
    wire N__10697;
    wire N__10696;
    wire N__10695;
    wire N__10694;
    wire N__10691;
    wire N__10690;
    wire N__10689;
    wire N__10688;
    wire N__10687;
    wire N__10686;
    wire N__10683;
    wire N__10682;
    wire N__10681;
    wire N__10680;
    wire N__10679;
    wire N__10676;
    wire N__10675;
    wire N__10674;
    wire N__10673;
    wire N__10672;
    wire N__10671;
    wire N__10670;
    wire N__10669;
    wire N__10668;
    wire N__10667;
    wire N__10666;
    wire N__10665;
    wire N__10664;
    wire N__10663;
    wire N__10662;
    wire N__10661;
    wire N__10658;
    wire N__10657;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10567;
    wire N__10564;
    wire N__10563;
    wire N__10562;
    wire N__10561;
    wire N__10560;
    wire N__10559;
    wire N__10558;
    wire N__10555;
    wire N__10554;
    wire N__10553;
    wire N__10552;
    wire N__10551;
    wire N__10550;
    wire N__10549;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10542;
    wire N__10535;
    wire N__10528;
    wire N__10525;
    wire N__10516;
    wire N__10511;
    wire N__10510;
    wire N__10509;
    wire N__10508;
    wire N__10507;
    wire N__10506;
    wire N__10505;
    wire N__10504;
    wire N__10501;
    wire N__10496;
    wire N__10493;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10489;
    wire N__10488;
    wire N__10487;
    wire N__10486;
    wire N__10481;
    wire N__10478;
    wire N__10471;
    wire N__10470;
    wire N__10469;
    wire N__10464;
    wire N__10453;
    wire N__10446;
    wire N__10439;
    wire N__10432;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10426;
    wire N__10425;
    wire N__10424;
    wire N__10417;
    wire N__10414;
    wire N__10413;
    wire N__10412;
    wire N__10409;
    wire N__10406;
    wire N__10395;
    wire N__10390;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10372;
    wire N__10369;
    wire N__10364;
    wire N__10359;
    wire N__10354;
    wire N__10351;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10270;
    wire N__10269;
    wire N__10268;
    wire N__10267;
    wire N__10266;
    wire N__10265;
    wire N__10264;
    wire N__10263;
    wire N__10262;
    wire N__10261;
    wire N__10260;
    wire N__10259;
    wire N__10258;
    wire N__10257;
    wire N__10256;
    wire N__10255;
    wire N__10254;
    wire N__10253;
    wire N__10252;
    wire N__10251;
    wire N__10250;
    wire N__10249;
    wire N__10248;
    wire N__10247;
    wire N__10246;
    wire N__10243;
    wire N__10242;
    wire N__10241;
    wire N__10240;
    wire N__10239;
    wire N__10238;
    wire N__10237;
    wire N__10236;
    wire N__10235;
    wire N__10234;
    wire N__10233;
    wire N__10232;
    wire N__10231;
    wire N__10230;
    wire N__10229;
    wire N__10228;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10113;
    wire N__10112;
    wire N__10107;
    wire N__10104;
    wire N__10101;
    wire N__10094;
    wire N__10091;
    wire N__10090;
    wire N__10089;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10079;
    wire N__10076;
    wire N__10071;
    wire N__10070;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10059;
    wire N__10056;
    wire N__10053;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10042;
    wire N__10041;
    wire N__10038;
    wire N__10035;
    wire N__10030;
    wire N__10029;
    wire N__10028;
    wire N__10025;
    wire N__10020;
    wire N__10017;
    wire N__10016;
    wire N__10013;
    wire N__10012;
    wire N__10011;
    wire N__10010;
    wire N__10007;
    wire N__10002;
    wire N__10001;
    wire N__10000;
    wire N__9999;
    wire N__9994;
    wire N__9993;
    wire N__9992;
    wire N__9989;
    wire N__9984;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9964;
    wire N__9959;
    wire N__9952;
    wire N__9949;
    wire N__9944;
    wire N__9937;
    wire N__9934;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9875;
    wire N__9872;
    wire N__9867;
    wire N__9864;
    wire N__9859;
    wire N__9858;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9846;
    wire N__9843;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9821;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9810;
    wire N__9809;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9768;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9749;
    wire N__9748;
    wire N__9747;
    wire N__9746;
    wire N__9741;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9713;
    wire N__9710;
    wire N__9709;
    wire N__9708;
    wire N__9705;
    wire N__9700;
    wire N__9699;
    wire N__9694;
    wire N__9691;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9655;
    wire N__9652;
    wire N__9651;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9638;
    wire N__9635;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9604;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9581;
    wire N__9572;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9560;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9529;
    wire N__9528;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9516;
    wire N__9513;
    wire N__9510;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9471;
    wire N__9468;
    wire N__9465;
    wire N__9462;
    wire N__9459;
    wire N__9456;
    wire N__9453;
    wire N__9450;
    wire N__9447;
    wire N__9444;
    wire N__9441;
    wire N__9436;
    wire N__9433;
    wire N__9428;
    wire N__9425;
    wire N__9422;
    wire N__9421;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9398;
    wire N__9395;
    wire N__9392;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9377;
    wire N__9374;
    wire N__9371;
    wire N__9370;
    wire N__9369;
    wire N__9366;
    wire N__9365;
    wire N__9364;
    wire N__9363;
    wire N__9356;
    wire N__9353;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9331;
    wire N__9328;
    wire N__9327;
    wire N__9326;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9285;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9242;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9226;
    wire N__9225;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9219;
    wire N__9218;
    wire N__9217;
    wire N__9216;
    wire N__9215;
    wire N__9214;
    wire N__9211;
    wire N__9210;
    wire N__9209;
    wire N__9206;
    wire N__9203;
    wire N__9200;
    wire N__9197;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9173;
    wire N__9170;
    wire N__9169;
    wire N__9168;
    wire N__9167;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9163;
    wire N__9162;
    wire N__9153;
    wire N__9152;
    wire N__9151;
    wire N__9150;
    wire N__9145;
    wire N__9138;
    wire N__9137;
    wire N__9134;
    wire N__9125;
    wire N__9116;
    wire N__9113;
    wire N__9106;
    wire N__9101;
    wire N__9098;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9064;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9056;
    wire N__9051;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9022;
    wire N__9017;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9009;
    wire N__9004;
    wire N__9001;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8968;
    wire N__8967;
    wire N__8964;
    wire N__8959;
    wire N__8956;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8872;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8857;
    wire N__8854;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8774;
    wire N__8771;
    wire N__8768;
    wire N__8767;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8725;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8702;
    wire N__8699;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8684;
    wire N__8681;
    wire N__8680;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8647;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8581;
    wire N__8580;
    wire N__8577;
    wire N__8572;
    wire N__8571;
    wire N__8570;
    wire N__8569;
    wire N__8564;
    wire N__8557;
    wire N__8552;
    wire N__8551;
    wire N__8550;
    wire N__8549;
    wire N__8548;
    wire N__8545;
    wire N__8542;
    wire N__8539;
    wire N__8536;
    wire N__8533;
    wire N__8522;
    wire N__8521;
    wire N__8520;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8512;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8493;
    wire N__8490;
    wire N__8485;
    wire N__8480;
    wire N__8473;
    wire N__8470;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8393;
    wire N__8390;
    wire N__8387;
    wire N__8384;
    wire N__8381;
    wire N__8378;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8350;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire N__8338;
    wire N__8337;
    wire N__8336;
    wire N__8333;
    wire N__8330;
    wire N__8329;
    wire N__8326;
    wire N__8323;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8303;
    wire N__8300;
    wire N__8299;
    wire N__8298;
    wire N__8297;
    wire N__8296;
    wire N__8295;
    wire N__8294;
    wire N__8291;
    wire N__8288;
    wire N__8285;
    wire N__8284;
    wire N__8281;
    wire N__8280;
    wire N__8277;
    wire N__8276;
    wire N__8275;
    wire N__8270;
    wire N__8267;
    wire N__8264;
    wire N__8261;
    wire N__8258;
    wire N__8253;
    wire N__8250;
    wire N__8245;
    wire N__8228;
    wire N__8227;
    wire N__8226;
    wire N__8225;
    wire N__8222;
    wire N__8221;
    wire N__8220;
    wire N__8217;
    wire N__8214;
    wire N__8213;
    wire N__8210;
    wire N__8207;
    wire N__8202;
    wire N__8197;
    wire N__8194;
    wire N__8183;
    wire N__8180;
    wire N__8177;
    wire N__8174;
    wire N__8171;
    wire N__8168;
    wire N__8165;
    wire N__8164;
    wire N__8161;
    wire N__8158;
    wire N__8153;
    wire N__8152;
    wire N__8151;
    wire N__8150;
    wire N__8149;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8139;
    wire N__8134;
    wire N__8131;
    wire N__8126;
    wire N__8125;
    wire N__8124;
    wire N__8121;
    wire N__8120;
    wire N__8119;
    wire N__8118;
    wire N__8117;
    wire N__8116;
    wire N__8115;
    wire N__8114;
    wire N__8113;
    wire N__8106;
    wire N__8101;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8082;
    wire N__8077;
    wire N__8074;
    wire N__8071;
    wire N__8054;
    wire N__8051;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8043;
    wire N__8042;
    wire N__8041;
    wire N__8040;
    wire N__8039;
    wire N__8038;
    wire N__8035;
    wire N__8034;
    wire N__8031;
    wire N__8026;
    wire N__8023;
    wire N__8022;
    wire N__8021;
    wire N__8020;
    wire N__8017;
    wire N__8016;
    wire N__8011;
    wire N__8008;
    wire N__8007;
    wire N__8006;
    wire N__8005;
    wire N__8004;
    wire N__8001;
    wire N__8000;
    wire N__7997;
    wire N__7992;
    wire N__7985;
    wire N__7984;
    wire N__7983;
    wire N__7982;
    wire N__7981;
    wire N__7980;
    wire N__7977;
    wire N__7974;
    wire N__7969;
    wire N__7960;
    wire N__7955;
    wire N__7948;
    wire N__7941;
    wire N__7936;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7906;
    wire N__7905;
    wire N__7902;
    wire N__7901;
    wire N__7898;
    wire N__7897;
    wire N__7894;
    wire N__7889;
    wire N__7888;
    wire N__7885;
    wire N__7880;
    wire N__7877;
    wire N__7876;
    wire N__7875;
    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7869;
    wire N__7866;
    wire N__7863;
    wire N__7860;
    wire N__7853;
    wire N__7848;
    wire N__7835;
    wire N__7832;
    wire N__7831;
    wire N__7828;
    wire N__7825;
    wire N__7820;
    wire N__7817;
    wire N__7816;
    wire N__7813;
    wire N__7810;
    wire N__7805;
    wire N__7802;
    wire N__7801;
    wire N__7798;
    wire N__7795;
    wire N__7790;
    wire N__7787;
    wire N__7786;
    wire N__7785;
    wire N__7784;
    wire N__7783;
    wire N__7782;
    wire N__7781;
    wire N__7772;
    wire N__7769;
    wire N__7764;
    wire N__7757;
    wire N__7754;
    wire N__7753;
    wire N__7750;
    wire N__7747;
    wire N__7744;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7732;
    wire N__7729;
    wire N__7726;
    wire N__7721;
    wire N__7718;
    wire N__7715;
    wire N__7712;
    wire N__7709;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7692;
    wire N__7687;
    wire N__7686;
    wire N__7685;
    wire N__7684;
    wire N__7683;
    wire N__7682;
    wire N__7679;
    wire N__7678;
    wire N__7677;
    wire N__7676;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7664;
    wire N__7659;
    wire N__7656;
    wire N__7651;
    wire N__7646;
    wire N__7631;
    wire N__7628;
    wire N__7627;
    wire N__7624;
    wire N__7623;
    wire N__7622;
    wire N__7619;
    wire N__7616;
    wire N__7613;
    wire N__7610;
    wire N__7601;
    wire N__7600;
    wire N__7599;
    wire N__7598;
    wire N__7593;
    wire N__7592;
    wire N__7591;
    wire N__7590;
    wire N__7589;
    wire N__7588;
    wire N__7587;
    wire N__7582;
    wire N__7581;
    wire N__7580;
    wire N__7577;
    wire N__7576;
    wire N__7575;
    wire N__7574;
    wire N__7571;
    wire N__7570;
    wire N__7569;
    wire N__7564;
    wire N__7559;
    wire N__7556;
    wire N__7553;
    wire N__7548;
    wire N__7545;
    wire N__7538;
    wire N__7531;
    wire N__7514;
    wire N__7511;
    wire N__7508;
    wire N__7505;
    wire N__7502;
    wire N__7499;
    wire N__7496;
    wire N__7493;
    wire N__7490;
    wire N__7489;
    wire N__7486;
    wire N__7485;
    wire N__7482;
    wire N__7479;
    wire N__7474;
    wire N__7469;
    wire N__7468;
    wire N__7467;
    wire N__7466;
    wire N__7463;
    wire N__7460;
    wire N__7457;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7443;
    wire N__7442;
    wire N__7439;
    wire N__7436;
    wire N__7433;
    wire N__7430;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7410;
    wire N__7407;
    wire N__7404;
    wire N__7401;
    wire N__7398;
    wire N__7395;
    wire N__7388;
    wire N__7385;
    wire N__7382;
    wire N__7379;
    wire N__7378;
    wire N__7377;
    wire N__7376;
    wire N__7375;
    wire N__7374;
    wire N__7371;
    wire N__7366;
    wire N__7363;
    wire N__7358;
    wire N__7349;
    wire N__7346;
    wire N__7343;
    wire N__7340;
    wire N__7337;
    wire N__7334;
    wire N__7333;
    wire N__7330;
    wire N__7329;
    wire N__7328;
    wire N__7325;
    wire N__7324;
    wire N__7323;
    wire N__7320;
    wire N__7317;
    wire N__7314;
    wire N__7309;
    wire N__7308;
    wire N__7307;
    wire N__7304;
    wire N__7299;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7287;
    wire N__7286;
    wire N__7285;
    wire N__7282;
    wire N__7277;
    wire N__7274;
    wire N__7265;
    wire N__7258;
    wire N__7247;
    wire N__7244;
    wire N__7241;
    wire N__7238;
    wire N__7235;
    wire N__7232;
    wire N__7229;
    wire N__7226;
    wire N__7223;
    wire N__7220;
    wire N__7217;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7190;
    wire N__7187;
    wire N__7184;
    wire N__7181;
    wire N__7178;
    wire N__7175;
    wire N__7172;
    wire N__7169;
    wire N__7166;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7130;
    wire N__7127;
    wire N__7124;
    wire N__7121;
    wire N__7118;
    wire N__7115;
    wire N__7112;
    wire N__7109;
    wire N__7106;
    wire N__7103;
    wire N__7100;
    wire N__7097;
    wire N__7094;
    wire N__7091;
    wire N__7088;
    wire N__7085;
    wire N__7082;
    wire N__7079;
    wire N__7076;
    wire N__7073;
    wire N__7070;
    wire N__7067;
    wire N__7064;
    wire N__7061;
    wire N__7060;
    wire N__7057;
    wire N__7054;
    wire N__7051;
    wire N__7048;
    wire N__7045;
    wire N__7040;
    wire N__7037;
    wire N__7036;
    wire N__7033;
    wire N__7032;
    wire N__7029;
    wire N__7026;
    wire N__7023;
    wire N__7020;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__7006;
    wire N__7003;
    wire N__6998;
    wire N__6997;
    wire N__6996;
    wire N__6993;
    wire N__6990;
    wire N__6987;
    wire N__6986;
    wire N__6985;
    wire N__6984;
    wire N__6981;
    wire N__6978;
    wire N__6975;
    wire N__6972;
    wire N__6969;
    wire N__6968;
    wire N__6967;
    wire N__6966;
    wire N__6963;
    wire N__6960;
    wire N__6953;
    wire N__6950;
    wire N__6945;
    wire N__6942;
    wire N__6929;
    wire N__6926;
    wire N__6923;
    wire N__6920;
    wire N__6917;
    wire N__6914;
    wire N__6911;
    wire N__6908;
    wire N__6905;
    wire N__6902;
    wire N__6901;
    wire N__6898;
    wire N__6897;
    wire N__6894;
    wire N__6891;
    wire N__6890;
    wire N__6889;
    wire N__6886;
    wire N__6883;
    wire N__6880;
    wire N__6877;
    wire N__6874;
    wire N__6871;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6845;
    wire N__6842;
    wire N__6839;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6827;
    wire N__6824;
    wire N__6821;
    wire N__6818;
    wire N__6815;
    wire N__6812;
    wire N__6809;
    wire N__6806;
    wire N__6803;
    wire N__6800;
    wire N__6797;
    wire N__6794;
    wire N__6791;
    wire N__6788;
    wire N__6785;
    wire N__6782;
    wire N__6779;
    wire N__6776;
    wire N__6773;
    wire N__6770;
    wire N__6767;
    wire N__6764;
    wire N__6761;
    wire N__6758;
    wire N__6755;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6730;
    wire N__6729;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6695;
    wire N__6694;
    wire N__6693;
    wire N__6690;
    wire N__6685;
    wire N__6680;
    wire N__6679;
    wire N__6676;
    wire N__6673;
    wire N__6668;
    wire N__6665;
    wire N__6662;
    wire N__6661;
    wire N__6656;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6619;
    wire N__6618;
    wire N__6615;
    wire N__6612;
    wire N__6609;
    wire N__6606;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6586;
    wire N__6581;
    wire N__6578;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6570;
    wire N__6565;
    wire N__6562;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6545;
    wire N__6542;
    wire N__6541;
    wire N__6540;
    wire N__6535;
    wire N__6532;
    wire N__6531;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6512;
    wire N__6509;
    wire N__6506;
    wire N__6503;
    wire N__6500;
    wire N__6499;
    wire N__6496;
    wire N__6493;
    wire N__6488;
    wire N__6485;
    wire N__6482;
    wire N__6479;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6471;
    wire N__6466;
    wire N__6461;
    wire N__6458;
    wire N__6457;
    wire N__6456;
    wire N__6455;
    wire N__6454;
    wire N__6451;
    wire N__6446;
    wire N__6443;
    wire N__6440;
    wire N__6431;
    wire N__6428;
    wire N__6425;
    wire N__6422;
    wire N__6421;
    wire N__6418;
    wire N__6415;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6391;
    wire N__6388;
    wire N__6385;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6364;
    wire N__6363;
    wire N__6360;
    wire N__6357;
    wire N__6354;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6325;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6312;
    wire N__6309;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6287;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6229;
    wire N__6226;
    wire N__6223;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6193;
    wire N__6190;
    wire N__6187;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6147;
    wire N__6142;
    wire N__6137;
    wire N__6134;
    wire N__6131;
    wire N__6128;
    wire N__6125;
    wire N__6124;
    wire N__6123;
    wire N__6120;
    wire N__6117;
    wire N__6114;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6100;
    wire N__6095;
    wire N__6094;
    wire N__6093;
    wire N__6090;
    wire N__6087;
    wire N__6084;
    wire N__6077;
    wire N__6076;
    wire N__6075;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6037;
    wire N__6034;
    wire N__6031;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6002;
    wire N__6001;
    wire N__5998;
    wire N__5995;
    wire N__5990;
    wire N__5987;
    wire N__5984;
    wire N__5981;
    wire N__5978;
    wire N__5975;
    wire N__5972;
    wire N__5971;
    wire N__5968;
    wire N__5965;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5953;
    wire N__5950;
    wire N__5947;
    wire N__5942;
    wire N__5941;
    wire N__5940;
    wire N__5939;
    wire N__5938;
    wire N__5937;
    wire N__5936;
    wire N__5931;
    wire N__5924;
    wire N__5919;
    wire N__5916;
    wire N__5909;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5897;
    wire N__5896;
    wire N__5893;
    wire N__5890;
    wire N__5885;
    wire N__5882;
    wire N__5881;
    wire N__5880;
    wire N__5875;
    wire N__5872;
    wire N__5871;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5855;
    wire N__5852;
    wire N__5849;
    wire N__5848;
    wire N__5847;
    wire N__5846;
    wire N__5845;
    wire N__5842;
    wire N__5841;
    wire N__5838;
    wire N__5837;
    wire N__5834;
    wire N__5827;
    wire N__5820;
    wire N__5819;
    wire N__5818;
    wire N__5815;
    wire N__5810;
    wire N__5805;
    wire N__5798;
    wire N__5797;
    wire N__5794;
    wire N__5791;
    wire N__5788;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5776;
    wire N__5773;
    wire N__5770;
    wire N__5765;
    wire N__5762;
    wire N__5759;
    wire N__5756;
    wire N__5753;
    wire N__5750;
    wire N__5747;
    wire N__5744;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5726;
    wire N__5723;
    wire N__5720;
    wire N__5717;
    wire N__5714;
    wire N__5711;
    wire N__5708;
    wire N__5705;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5684;
    wire N__5681;
    wire N__5678;
    wire N__5675;
    wire N__5672;
    wire N__5671;
    wire N__5670;
    wire N__5669;
    wire N__5668;
    wire N__5667;
    wire N__5664;
    wire N__5661;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5636;
    wire N__5633;
    wire N__5626;
    wire N__5621;
    wire N__5618;
    wire N__5615;
    wire N__5612;
    wire N__5609;
    wire N__5606;
    wire N__5603;
    wire N__5602;
    wire N__5599;
    wire N__5596;
    wire N__5591;
    wire N__5588;
    wire N__5585;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5524;
    wire N__5523;
    wire N__5520;
    wire N__5515;
    wire N__5510;
    wire N__5509;
    wire N__5508;
    wire N__5505;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5491;
    wire N__5488;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5468;
    wire N__5465;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5450;
    wire N__5447;
    wire N__5446;
    wire N__5443;
    wire N__5440;
    wire N__5435;
    wire N__5434;
    wire N__5431;
    wire N__5428;
    wire N__5425;
    wire N__5422;
    wire N__5419;
    wire N__5416;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5404;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5339;
    wire N__5336;
    wire N__5333;
    wire N__5330;
    wire N__5327;
    wire N__5324;
    wire N__5321;
    wire N__5318;
    wire N__5317;
    wire N__5314;
    wire N__5311;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5299;
    wire N__5296;
    wire N__5293;
    wire N__5290;
    wire N__5287;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5275;
    wire N__5270;
    wire N__5267;
    wire N__5266;
    wire N__5265;
    wire N__5262;
    wire N__5257;
    wire N__5252;
    wire N__5249;
    wire N__5248;
    wire N__5245;
    wire N__5242;
    wire N__5241;
    wire N__5238;
    wire N__5235;
    wire N__5232;
    wire N__5229;
    wire N__5226;
    wire N__5223;
    wire N__5220;
    wire N__5217;
    wire N__5214;
    wire N__5209;
    wire N__5206;
    wire N__5205;
    wire N__5200;
    wire N__5197;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5162;
    wire N__5159;
    wire N__5156;
    wire N__5155;
    wire N__5152;
    wire N__5149;
    wire N__5144;
    wire N__5143;
    wire N__5142;
    wire N__5141;
    wire N__5136;
    wire N__5131;
    wire N__5126;
    wire N__5123;
    wire N__5120;
    wire N__5117;
    wire N__5116;
    wire N__5115;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5066;
    wire N__5063;
    wire N__5060;
    wire N__5059;
    wire N__5056;
    wire N__5053;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5011;
    wire N__5008;
    wire N__5005;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4973;
    wire N__4970;
    wire N__4967;
    wire N__4964;
    wire N__4961;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4933;
    wire N__4932;
    wire N__4929;
    wire N__4924;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4895;
    wire N__4892;
    wire N__4891;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4852;
    wire N__4849;
    wire N__4846;
    wire N__4843;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4819;
    wire N__4816;
    wire N__4815;
    wire N__4810;
    wire N__4807;
    wire N__4802;
    wire N__4801;
    wire N__4798;
    wire N__4795;
    wire N__4792;
    wire N__4787;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4760;
    wire N__4757;
    wire N__4754;
    wire N__4753;
    wire N__4750;
    wire N__4747;
    wire N__4742;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4730;
    wire N__4727;
    wire N__4724;
    wire N__4721;
    wire N__4718;
    wire N__4717;
    wire N__4714;
    wire N__4711;
    wire N__4708;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4694;
    wire N__4691;
    wire N__4688;
    wire N__4685;
    wire N__4682;
    wire N__4679;
    wire N__4676;
    wire N__4673;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4655;
    wire N__4652;
    wire N__4649;
    wire N__4646;
    wire N__4643;
    wire N__4640;
    wire N__4637;
    wire N__4634;
    wire N__4631;
    wire N__4628;
    wire N__4625;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4600;
    wire N__4599;
    wire N__4598;
    wire N__4597;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4579;
    wire N__4576;
    wire N__4573;
    wire N__4568;
    wire N__4567;
    wire N__4564;
    wire N__4561;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4486;
    wire N__4483;
    wire N__4480;
    wire N__4477;
    wire N__4474;
    wire N__4471;
    wire N__4468;
    wire N__4465;
    wire N__4462;
    wire N__4461;
    wire N__4458;
    wire N__4455;
    wire N__4452;
    wire N__4447;
    wire N__4444;
    wire N__4443;
    wire N__4438;
    wire N__4435;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire CLK40_IN_c;
    wire VCCG0;
    wire GNDG0;
    wire CLK80_PLL_i_i;
    wire DBRn_c_i_0;
    wire VBENn_c;
    wire A_c_14;
    wire CMA_c_1;
    wire \U712_CHIP_RAM.N_340 ;
    wire CMA_c_5;
    wire \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ;
    wire \U712_CHIP_RAM.N_297_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ;
    wire \U712_CHIP_RAM.N_196_cascade_ ;
    wire TACK_EN;
    wire \U712_CHIP_RAM.REFRESH5lto0 ;
    wire bfn_9_5_0_;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ;
    wire C1_c_g;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ;
    wire A_c_16;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ;
    wire A_c_10;
    wire \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ;
    wire CMA_c_7;
    wire CMA_c_8;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0 ;
    wire \U712_CHIP_RAM.N_556_cascade_ ;
    wire \U712_CHIP_RAM.N_202 ;
    wire \U712_CHIP_RAM.N_388_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0 ;
    wire \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.REFRESH5lto7_0 ;
    wire \U712_CHIP_RAM.REFRESH5lt7 ;
    wire \U712_CHIP_RAM.REFRESHZ0 ;
    wire RAMSPACEn_c;
    wire \U712_CHIP_RAM.N_417_cascade_ ;
    wire \U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ;
    wire \U712_CHIP_RAM.N_206 ;
    wire \U712_CHIP_RAM.N_457 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_5 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_4 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1 ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ;
    wire LATCH_CLK_c;
    wire TSn_c;
    wire REGSPACEn_c;
    wire \U712_REG_SM.N_414 ;
    wire \U712_CYCLE_TERM.N_452_cascade_ ;
    wire \U712_CYCLE_TERM.N_312 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ1Z_2 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_3 ;
    wire TACK_OUTn;
    wire DBRn_c;
    wire DBR_SYNCZ0Z_0;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_4 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_1 ;
    wire \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ;
    wire \U712_CYCLE_TERM.TACK_STATEZ0Z_0 ;
    wire C3_c;
    wire \U712_REG_SM.START_RSTZ0 ;
    wire C1_c;
    wire \U712_REG_SM.C1_SYNCZ0Z_0 ;
    wire CRCSn_c;
    wire RASn_c;
    wire CMA_c_0;
    wire CMA_c_10;
    wire CMA_c_2;
    wire A_c_9;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ;
    wire A_c_17;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ;
    wire \U712_CHIP_RAM.N_346 ;
    wire \U712_CHIP_RAM.N_388 ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ;
    wire \U712_CHIP_RAM.REFRESH_RST ;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ;
    wire \U712_CHIP_RAM.N_445 ;
    wire \U712_CHIP_RAM.N_208 ;
    wire \U712_CHIP_RAM.N_303 ;
    wire \U712_CHIP_RAM.N_443_cascade_ ;
    wire \U712_CHIP_RAM.N_204 ;
    wire \U712_CHIP_RAM.N_463_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ;
    wire \U712_CHIP_RAM.N_439 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ;
    wire CLK_EN_c;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ;
    wire \U712_CHIP_RAM.N_360 ;
    wire \U712_CHIP_RAM.N_418 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0 ;
    wire \U712_REG_SM.N_400_cascade_ ;
    wire \U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ;
    wire \U712_CHIP_RAM.N_405 ;
    wire bfn_10_12_0_;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ;
    wire \U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ;
    wire CPU_TACKm;
    wire \U712_CYCLE_TERM.TACK_EN6_0 ;
    wire DBR_SYNCZ0Z_1;
    wire DBR_SYNC_i_1;
    wire \U712_REG_SM.N_307_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_3 ;
    wire REGENn_c;
    wire \U712_REG_SM.REGENn_e_1 ;
    wire \U712_REG_SM.REG_CYCLE_STARTZ0 ;
    wire \U712_REG_SM.WRITE_CYCLEZ0 ;
    wire A_c_12;
    wire A_c_11;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ;
    wire \U712_CHIP_RAM.N_551 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ;
    wire A_c_20;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.N_555_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER16 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ;
    wire \U712_CHIP_RAM.N_556 ;
    wire \U712_CHIP_RAM.N_302 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER19 ;
    wire \U712_CHIP_RAM.N_355_cascade_ ;
    wire \U712_CHIP_RAM.N_389 ;
    wire \U712_CHIP_RAM.N_301 ;
    wire \U712_CHIP_RAM.N_289 ;
    wire \U712_CHIP_RAM.N_356 ;
    wire \U712_CHIP_RAM.N_356_cascade_ ;
    wire \U712_CHIP_RAM.N_448 ;
    wire \U712_CHIP_RAM.N_288_cascade_ ;
    wire \U712_CHIP_RAM.N_473 ;
    wire \U712_CHIP_RAM.N_473_cascade_ ;
    wire \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0 ;
    wire \U712_CHIP_RAM.N_362 ;
    wire \U712_CHIP_RAM.N_463 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ;
    wire \U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ;
    wire DBDIR_c;
    wire \U712_CHIP_RAM.CAS_SYNCZ0Z_0 ;
    wire \U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ;
    wire \U712_REG_SM.N_306_cascade_ ;
    wire \U712_REG_SM.N_399_cascade_ ;
    wire \U712_REG_SM.REG_CYCLE_5_iv_0_0 ;
    wire \U712_REG_SM.N_311 ;
    wire \U712_REG_SM.N_353_cascade_ ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_2 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_0 ;
    wire \U712_REG_SM.N_322 ;
    wire REG_TACK;
    wire \U712_REG_SM.STATE_COUNTsr_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_0 ;
    wire \U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_7 ;
    wire \U712_REG_SM.N_307 ;
    wire \U712_REG_SM.N_553 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_4 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_5 ;
    wire \U712_REG_SM.STATE_COUNTZ1Z_6 ;
    wire N_130_i;
    wire CONSTANT_ONE_NET;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ;
    wire WEn_c;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ;
    wire A_c_13;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ;
    wire A_c_15;
    wire \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ;
    wire A_c_6;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ;
    wire A_c_2;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ;
    wire A_c_3;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ;
    wire A_c_4;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ;
    wire A_c_7;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ;
    wire A_c_8;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ;
    wire A_c_18;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ;
    wire A_c_5;
    wire \U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ;
    wire AWEn_c;
    wire \U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ;
    wire \U712_CHIP_RAM.N_294_cascade_ ;
    wire \U712_CHIP_RAM.N_288 ;
    wire \U712_CHIP_RAM.N_469_cascade_ ;
    wire \U712_CHIP_RAM.N_557 ;
    wire \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ;
    wire \U712_CHIP_RAM.N_555 ;
    wire \U712_CHIP_RAM.N_309_cascade_ ;
    wire \U712_CHIP_RAM.N_387 ;
    wire \U712_CHIP_RAM.N_200_cascade_ ;
    wire \U712_CHIP_RAM.N_309 ;
    wire \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ;
    wire \U712_CHIP_RAM.WRITE_CYCLEZ0 ;
    wire \U712_CHIP_RAM.N_285 ;
    wire \U712_CHIP_RAM.N_285_cascade_ ;
    wire \U712_CHIP_RAM.N_293 ;
    wire \U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_0 ;
    wire bfn_12_9_0_;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_s_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ;
    wire \U712_CHIP_RAM.N_200 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ;
    wire \U712_CHIP_RAM.SDRAM_COUNTERe_0_i ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_3 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_1 ;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_2 ;
    wire \U712_BYTE_ENABLE.N_451 ;
    wire N_211_i;
    wire \U712_BYTE_ENABLE.N_410_cascade_ ;
    wire N_148_i;
    wire \U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_1 ;
    wire \U712_REG_SM.C3_SYNCZ0Z_1 ;
    wire \U712_REG_SM.STATE_COUNTZ0Z_8 ;
    wire \U712_REG_SM.N_95_cascade_ ;
    wire \U712_REG_SM.N_432 ;
    wire LDSn_c;
    wire \U712_REG_SM.N_95 ;
    wire UDSn_c;
    wire \U712_REG_SM.N_433 ;
    wire RESETn_c_i;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ;
    wire CMA_c_3;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ;
    wire CMA_c_4;
    wire \U712_CHIP_RAM.N_297 ;
    wire \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ;
    wire \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ;
    wire CMA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_AZ0Z1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ;
    wire \INVU712_CHIP_RAM.DMA_A1_nesrC_net ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ;
    wire DBRn_c_i;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ;
    wire \U712_BYTE_ENABLE.N_409 ;
    wire \U712_REG_SM.C1_SYNCZ0Z_1 ;
    wire ASn_c;
    wire \U712_REG_SM.N_95_0 ;
    wire LLBEn_c;
    wire \U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ;
    wire CASn_c;
    wire DRA_c_5;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ;
    wire DRA_c_2;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ;
    wire DRA_c_1;
    wire DRA_c_0;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ;
    wire DRA_c_8;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ;
    wire DRA_c_7;
    wire DRA_c_6;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ;
    wire \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ;
    wire \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ;
    wire DRA_c_4;
    wire DRA_c_3;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ;
    wire N_146_i;
    wire CLK40_PLL_i;
    wire CLK40_PLL_i_i;
    wire \U712_BYTE_ENABLE.N_406 ;
    wire \U712_BYTE_ENABLE.N_284_i ;
    wire N_374_i;
    wire N_373_i;
    wire A_c_1;
    wire A_c_0;
    wire SIZ_c_0;
    wire SIZ_c_1;
    wire UMBEn_c;
    wire \U712_CHIP_RAM.CMA_5_i_0_9 ;
    wire A_c_19;
    wire CMA_c_9;
    wire \U712_CHIP_RAM.un1_CMA25_0_i_0 ;
    wire DMA_CYCLEm;
    wire \U712_BYTE_ENABLE.N_411 ;
    wire DBENn_c;
    wire N_150_i;
    wire AGNUS_REV_c;
    wire DRA_c_9;
    wire \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ;
    wire C3_c_g;
    wire DBRn_c_i_0_g;
    wire RESETn_c_i_g;
    wire RESETn_c;
    wire RAS1n_c;
    wire RAS0n_c;
    wire \U712_CHIP_RAM.RAS_SYNCZ0Z_0 ;
    wire CLK80_PLL;
    wire REG_CYCLEm;
    wire CPU_CYCLEm;
    wire N_136_i;
    wire CASUn_c;
    wire RnW_c;
    wire CASLn_c;
    wire DMA_WRITE_CYCLE;
    wire N_357;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam pll.PLLOUT_SELECT_PORTA="GENCLK";
    defparam pll.FILTER_RANGE=3'b011;
    defparam pll.FEEDBACK_PATH="DELAY";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE_PORTB=1'b0;
    defparam pll.ENABLE_ICEGATE_PORTA=1'b0;
    defparam pll.DIVR=4'b0000;
    defparam pll.DIVQ=3'b011;
    defparam pll.DIVF=7'b0000001;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE pll (
            .EXTFEEDBACK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(CLK40_PLL_i),
            .REFERENCECLK(N__4376),
            .RESETB(N__6917),
            .BYPASS(),
            .PLLOUTCOREA(),
            .SDI(),
            .PLLOUTGLOBALB(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(),
            .PLLOUTGLOBALA(CLK80_PLL),
            .SCLK());
    IO_PAD DBENn_obuf_iopad (
            .OE(N__12615),
            .DIN(N__12614),
            .DOUT(N__12613),
            .PACKAGEPIN(DBENn));
    defparam DBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBENn_obuf_preio (
            .PADOEN(N__12615),
            .PADOUT(N__12614),
            .PADIN(N__12613),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11093),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_2_iopad (
            .OE(N__12606),
            .DIN(N__12605),
            .DOUT(N__12604),
            .PACKAGEPIN(A[2]));
    defparam A_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_2_preio (
            .PADOEN(N__12606),
            .PADOUT(N__12605),
            .PADIN(N__12604),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASn_obuf_iopad (
            .OE(N__12597),
            .DIN(N__12596),
            .DOUT(N__12595),
            .PACKAGEPIN(CASn));
    defparam CASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CASn_obuf_preio (
            .PADOEN(N__12597),
            .PADOUT(N__12596),
            .PADIN(N__12595),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9083),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDDIR_obuf_iopad (
            .OE(N__12588),
            .DIN(N__12587),
            .DOUT(N__12586),
            .PACKAGEPIN(DRDDIR));
    defparam DRDDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDDIR_obuf_preio (
            .PADOEN(N__12588),
            .PADOUT(N__12587),
            .PADIN(N__12586),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11651),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C1_ibuf_iopad (
            .OE(N__12579),
            .DIN(N__12578),
            .DOUT(N__12577),
            .PACKAGEPIN(C1));
    defparam C1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C1_ibuf_preio (
            .PADOEN(N__12579),
            .PADOUT(N__12578),
            .PADIN(N__12577),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK1_obuf_iopad (
            .OE(N__12570),
            .DIN(N__12569),
            .DOUT(N__12568),
            .PACKAGEPIN(BANK1));
    defparam BANK1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK1_obuf_preio (
            .PADOEN(N__12570),
            .PADOUT(N__12569),
            .PADIN(N__12568),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_3_iopad (
            .OE(N__12561),
            .DIN(N__12560),
            .DOUT(N__12559),
            .PACKAGEPIN(DRA[3]));
    defparam DRA_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_3_preio (
            .PADOEN(N__12561),
            .PADOUT(N__12560),
            .PADIN(N__12559),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AGNUS_REV_ibuf_iopad (
            .OE(N__12552),
            .DIN(N__12551),
            .DOUT(N__12550),
            .PACKAGEPIN(AGNUS_REV));
    defparam AGNUS_REV_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AGNUS_REV_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AGNUS_REV_ibuf_preio (
            .PADOEN(N__12552),
            .PADOUT(N__12551),
            .PADIN(N__12550),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AGNUS_REV_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS0n_ibuf_iopad (
            .OE(N__12543),
            .DIN(N__12542),
            .DOUT(N__12541),
            .PACKAGEPIN(RAS0n));
    defparam RAS0n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS0n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS0n_ibuf_preio (
            .PADOEN(N__12543),
            .PADOUT(N__12542),
            .PADIN(N__12541),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS0n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAS1n_ibuf_iopad (
            .OE(N__12534),
            .DIN(N__12533),
            .DOUT(N__12532),
            .PACKAGEPIN(RAS1n));
    defparam RAS1n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAS1n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAS1n_ibuf_preio (
            .PADOEN(N__12534),
            .PADOUT(N__12533),
            .PADIN(N__12532),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAS1n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_7_iopad (
            .OE(N__12525),
            .DIN(N__12524),
            .DOUT(N__12523),
            .PACKAGEPIN(A[7]));
    defparam A_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_7_preio (
            .PADOEN(N__12525),
            .PADOUT(N__12524),
            .PADIN(N__12523),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_7_iopad (
            .OE(N__12516),
            .DIN(N__12515),
            .DOUT(N__12514),
            .PACKAGEPIN(CMA[7]));
    defparam CMA_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_7_preio (
            .PADOEN(N__12516),
            .PADOUT(N__12515),
            .PADIN(N__12514),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4673),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UUBEn_obuf_iopad (
            .OE(N__12507),
            .DIN(N__12506),
            .DOUT(N__12505),
            .PACKAGEPIN(UUBEn));
    defparam UUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UUBEn_obuf_preio (
            .PADOEN(N__12507),
            .PADOUT(N__12506),
            .PADIN(N__12505),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11633),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_9_iopad (
            .OE(N__12498),
            .DIN(N__12497),
            .DOUT(N__12496),
            .PACKAGEPIN(DRA[9]));
    defparam DRA_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_9_preio (
            .PADOEN(N__12498),
            .PADOUT(N__12497),
            .PADIN(N__12496),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGSPACEn_ibuf_iopad (
            .OE(N__12489),
            .DIN(N__12488),
            .DOUT(N__12487),
            .PACKAGEPIN(REGSPACEn));
    defparam REGSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam REGSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO REGSPACEn_ibuf_preio (
            .PADOEN(N__12489),
            .PADOUT(N__12488),
            .PADIN(N__12487),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(REGSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_0_iopad (
            .OE(N__12480),
            .DIN(N__12479),
            .DOUT(N__12478),
            .PACKAGEPIN(SIZ[0]));
    defparam SIZ_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_0_preio (
            .PADOEN(N__12480),
            .PADOUT(N__12479),
            .PADIN(N__12478),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VBENn_obuf_iopad (
            .OE(N__12471),
            .DIN(N__12470),
            .DOUT(N__12469),
            .PACKAGEPIN(VBENn));
    defparam VBENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VBENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VBENn_obuf_preio (
            .PADOEN(N__12471),
            .PADOUT(N__12470),
            .PADIN(N__12469),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4406),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASUn_ibuf_iopad (
            .OE(N__12462),
            .DIN(N__12461),
            .DOUT(N__12460),
            .PACKAGEPIN(CASUn));
    defparam CASUn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASUn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASUn_ibuf_preio (
            .PADOEN(N__12462),
            .PADOUT(N__12461),
            .PADIN(N__12460),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASUn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_4_iopad (
            .OE(N__12453),
            .DIN(N__12452),
            .DOUT(N__12451),
            .PACKAGEPIN(A[4]));
    defparam A_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_4_preio (
            .PADOEN(N__12453),
            .PADOUT(N__12452),
            .PADIN(N__12451),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_0_iopad (
            .OE(N__12444),
            .DIN(N__12443),
            .DOUT(N__12442),
            .PACKAGEPIN(CMA[0]));
    defparam CMA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_0_preio (
            .PADOEN(N__12444),
            .PADOUT(N__12443),
            .PADIN(N__12442),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5354),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBRn_ibuf_iopad (
            .OE(N__12435),
            .DIN(N__12434),
            .DOUT(N__12433),
            .PACKAGEPIN(DBRn));
    defparam DBRn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam DBRn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO DBRn_ibuf_preio (
            .PADOEN(N__12435),
            .PADOUT(N__12434),
            .PADIN(N__12433),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DBRn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CRCSn_obuf_iopad (
            .OE(N__12426),
            .DIN(N__12425),
            .DOUT(N__12424),
            .PACKAGEPIN(CRCSn));
    defparam CRCSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CRCSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CRCSn_obuf_preio (
            .PADOEN(N__12426),
            .PADOUT(N__12425),
            .PADIN(N__12424),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5393),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_12_iopad (
            .OE(N__12417),
            .DIN(N__12416),
            .DOUT(N__12415),
            .PACKAGEPIN(A[12]));
    defparam A_ibuf_12_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_12_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_12_preio (
            .PADOEN(N__12417),
            .PADOUT(N__12416),
            .PADIN(N__12415),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_12),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LLBEn_obuf_iopad (
            .OE(N__12408),
            .DIN(N__12407),
            .DOUT(N__12406),
            .PACKAGEPIN(LLBEn));
    defparam LLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LLBEn_obuf_preio (
            .PADOEN(N__12408),
            .PADOUT(N__12407),
            .PADIN(N__12406),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9242),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TBIn_obuft_iopad (
            .OE(N__12399),
            .DIN(N__12398),
            .DOUT(N__12397),
            .PACKAGEPIN(TBIn));
    defparam TBIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TBIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TBIn_obuft_preio (
            .PADOEN(N__12399),
            .PADOUT(N__12398),
            .PADIN(N__12397),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4486),
            .DIN0(),
            .DOUT0(N__5248),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CASLn_ibuf_iopad (
            .OE(N__12390),
            .DIN(N__12389),
            .DOUT(N__12388),
            .PACKAGEPIN(CASLn));
    defparam CASLn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CASLn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CASLn_ibuf_preio (
            .PADOEN(N__12390),
            .PADOUT(N__12389),
            .PADIN(N__12388),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CASLn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TSn_ibuf_iopad (
            .OE(N__12381),
            .DIN(N__12380),
            .DOUT(N__12379),
            .PACKAGEPIN(TSn));
    defparam TSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam TSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO TSn_ibuf_preio (
            .PADOEN(N__12381),
            .PADOUT(N__12380),
            .PADIN(N__12379),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TSn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RAMSPACEn_ibuf_iopad (
            .OE(N__12372),
            .DIN(N__12371),
            .DOUT(N__12370),
            .PACKAGEPIN(RAMSPACEn));
    defparam RAMSPACEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RAMSPACEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RAMSPACEn_ibuf_preio (
            .PADOEN(N__12372),
            .PADOUT(N__12371),
            .PADIN(N__12370),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RAMSPACEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_18_iopad (
            .OE(N__12363),
            .DIN(N__12362),
            .DOUT(N__12361),
            .PACKAGEPIN(A[18]));
    defparam A_ibuf_18_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_18_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_18_preio (
            .PADOEN(N__12363),
            .PADOUT(N__12362),
            .PADIN(N__12361),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_18),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_9_iopad (
            .OE(N__12354),
            .DIN(N__12353),
            .DOUT(N__12352),
            .PACKAGEPIN(A[9]));
    defparam A_ibuf_9_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_9_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_9_preio (
            .PADOEN(N__12354),
            .PADOUT(N__12353),
            .PADIN(N__12352),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DMA_LATCH_EN_obuf_iopad (
            .OE(N__12345),
            .DIN(N__12344),
            .DOUT(N__12343),
            .PACKAGEPIN(DMA_LATCH_EN));
    defparam DMA_LATCH_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DMA_LATCH_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DMA_LATCH_EN_obuf_preio (
            .PADOEN(N__12345),
            .PADOUT(N__12344),
            .PADIN(N__12343),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6647),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_7_iopad (
            .OE(N__12336),
            .DIN(N__12335),
            .DOUT(N__12334),
            .PACKAGEPIN(DRA[7]));
    defparam DRA_ibuf_7_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_7_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_7_preio (
            .PADOEN(N__12336),
            .PADOUT(N__12335),
            .PADIN(N__12334),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_15_iopad (
            .OE(N__12327),
            .DIN(N__12326),
            .DOUT(N__12325),
            .PACKAGEPIN(A[15]));
    defparam A_ibuf_15_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_15_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_15_preio (
            .PADOEN(N__12327),
            .PADOUT(N__12326),
            .PADIN(N__12325),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_15),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RESETn_ibuf_iopad (
            .OE(N__12318),
            .DIN(N__12317),
            .DOUT(N__12316),
            .PACKAGEPIN(RESETn));
    defparam RESETn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RESETn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RESETn_ibuf_preio (
            .PADOEN(N__12318),
            .PADOUT(N__12317),
            .PADIN(N__12316),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RESETn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_3_iopad (
            .OE(N__12309),
            .DIN(N__12308),
            .DOUT(N__12307),
            .PACKAGEPIN(A[3]));
    defparam A_ibuf_3_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_3_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_3_preio (
            .PADOEN(N__12309),
            .PADOUT(N__12308),
            .PADIN(N__12307),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40_IN_ibuf_iopad (
            .OE(N__12300),
            .DIN(N__12299),
            .DOUT(N__12298),
            .PACKAGEPIN(CLK40_IN));
    defparam CLK40_IN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40_IN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK40_IN_ibuf_preio (
            .PADOEN(N__12300),
            .PADOUT(N__12299),
            .PADIN(N__12298),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(CLK40_IN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RASn_obuf_iopad (
            .OE(N__12291),
            .DIN(N__12290),
            .DOUT(N__12289),
            .PACKAGEPIN(RASn));
    defparam RASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RASn_obuf_preio (
            .PADOEN(N__12291),
            .PADOUT(N__12290),
            .PADIN(N__12289),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5372),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BANK0_obuf_iopad (
            .OE(N__12282),
            .DIN(N__12281),
            .DOUT(N__12280),
            .PACKAGEPIN(BANK0));
    defparam BANK0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam BANK0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO BANK0_obuf_preio (
            .PADOEN(N__12282),
            .PADOUT(N__12281),
            .PADIN(N__12280),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_0_iopad (
            .OE(N__12273),
            .DIN(N__12272),
            .DOUT(N__12271),
            .PACKAGEPIN(DRA[0]));
    defparam DRA_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_0_preio (
            .PADOEN(N__12273),
            .PADOUT(N__12272),
            .PADIN(N__12271),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD ASn_obuf_iopad (
            .OE(N__12264),
            .DIN(N__12263),
            .DOUT(N__12262),
            .PACKAGEPIN(ASn));
    defparam ASn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam ASn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO ASn_obuf_preio (
            .PADOEN(N__12264),
            .PADOUT(N__12263),
            .PADIN(N__12262),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9266),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_0_iopad (
            .OE(N__12255),
            .DIN(N__12254),
            .DOUT(N__12253),
            .PACKAGEPIN(DA[0]));
    defparam DA_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_0_preio (
            .PADOEN(N__12255),
            .PADOUT(N__12254),
            .PADIN(N__12253),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5318),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_0_iopad (
            .OE(N__12246),
            .DIN(N__12245),
            .DOUT(N__12244),
            .PACKAGEPIN(A[0]));
    defparam A_ibuf_0_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_0_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_0_preio (
            .PADOEN(N__12246),
            .PADOUT(N__12245),
            .PADIN(N__12244),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_0),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_10_iopad (
            .OE(N__12237),
            .DIN(N__12236),
            .DOUT(N__12235),
            .PACKAGEPIN(CMA[10]));
    defparam CMA_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_10_preio (
            .PADOEN(N__12237),
            .PADOUT(N__12236),
            .PADIN(N__12235),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5342),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_4_iopad (
            .OE(N__12228),
            .DIN(N__12227),
            .DOUT(N__12226),
            .PACKAGEPIN(CMA[4]));
    defparam CMA_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_4_preio (
            .PADOEN(N__12228),
            .PADOUT(N__12227),
            .PADIN(N__12226),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD REGENn_obuf_iopad (
            .OE(N__12219),
            .DIN(N__12218),
            .DOUT(N__12217),
            .PACKAGEPIN(REGENn));
    defparam REGENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam REGENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO REGENn_obuf_preio (
            .PADOEN(N__12219),
            .PADOUT(N__12218),
            .PADIN(N__12217),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6137),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_19_iopad (
            .OE(N__12210),
            .DIN(N__12209),
            .DOUT(N__12208),
            .PACKAGEPIN(A[19]));
    defparam A_ibuf_19_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_19_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_19_preio (
            .PADOEN(N__12210),
            .PADOUT(N__12209),
            .PADIN(N__12208),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_19),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_8_iopad (
            .OE(N__12201),
            .DIN(N__12200),
            .DOUT(N__12199),
            .PACKAGEPIN(A[8]));
    defparam A_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_8_preio (
            .PADOEN(N__12201),
            .PADOUT(N__12200),
            .PADIN(N__12199),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLMBEn_obuf_iopad (
            .OE(N__12192),
            .DIN(N__12191),
            .DOUT(N__12190),
            .PACKAGEPIN(CLMBEn));
    defparam CLMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLMBEn_obuf_preio (
            .PADOEN(N__12192),
            .PADOUT(N__12191),
            .PADIN(N__12190),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11021),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TCIn_obuft_iopad (
            .OE(N__12183),
            .DIN(N__12182),
            .DOUT(N__12181),
            .PACKAGEPIN(TCIn));
    defparam TCIn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TCIn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TCIn_obuft_preio (
            .PADOEN(N__12183),
            .PADOUT(N__12182),
            .PADIN(N__12181),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4487),
            .DIN0(),
            .DOUT0(N__5252),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD WEn_obuf_iopad (
            .OE(N__12174),
            .DIN(N__12173),
            .DOUT(N__12172),
            .PACKAGEPIN(WEn));
    defparam WEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam WEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO WEn_obuf_preio (
            .PADOEN(N__12174),
            .PADOUT(N__12173),
            .PADIN(N__12172),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6860),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DBDIR_obuf_iopad (
            .OE(N__12165),
            .DIN(N__12164),
            .DOUT(N__12163),
            .PACKAGEPIN(DBDIR));
    defparam DBDIR_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DBDIR_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DBDIR_obuf_preio (
            .PADOEN(N__12165),
            .PADOUT(N__12164),
            .PADIN(N__12163),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6407),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUMBEn_obuf_iopad (
            .OE(N__12156),
            .DIN(N__12155),
            .DOUT(N__12154),
            .PACKAGEPIN(CUMBEn));
    defparam CUMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUMBEn_obuf_preio (
            .PADOEN(N__12156),
            .PADOUT(N__12155),
            .PADIN(N__12154),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8369),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_6_iopad (
            .OE(N__12147),
            .DIN(N__12146),
            .DOUT(N__12145),
            .PACKAGEPIN(DRA[6]));
    defparam DRA_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_6_preio (
            .PADOEN(N__12147),
            .PADOUT(N__12146),
            .PADIN(N__12145),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_5_iopad (
            .OE(N__12138),
            .DIN(N__12137),
            .DOUT(N__12136),
            .PACKAGEPIN(A[5]));
    defparam A_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_5_preio (
            .PADOEN(N__12138),
            .PADOUT(N__12137),
            .PADIN(N__12136),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_2_iopad (
            .OE(N__12129),
            .DIN(N__12128),
            .DOUT(N__12127),
            .PACKAGEPIN(DA[2]));
    defparam DA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_2_preio (
            .PADOEN(N__12129),
            .PADOUT(N__12128),
            .PADIN(N__12127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6047),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RnW_ibuf_iopad (
            .OE(N__12120),
            .DIN(N__12119),
            .DOUT(N__12118),
            .PACKAGEPIN(RnW));
    defparam RnW_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam RnW_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO RnW_ibuf_preio (
            .PADOEN(N__12120),
            .PADOUT(N__12119),
            .PADIN(N__12118),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(RnW_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_16_iopad (
            .OE(N__12111),
            .DIN(N__12110),
            .DOUT(N__12109),
            .PACKAGEPIN(A[16]));
    defparam A_ibuf_16_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_16_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_16_preio (
            .PADOEN(N__12111),
            .PADOUT(N__12110),
            .PADIN(N__12109),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_16),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_1_iopad (
            .OE(N__12102),
            .DIN(N__12101),
            .DOUT(N__12100),
            .PACKAGEPIN(CMA[1]));
    defparam CMA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_1_preio (
            .PADOEN(N__12102),
            .PADOUT(N__12101),
            .PADIN(N__12100),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4556),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LMBEn_obuf_iopad (
            .OE(N__12093),
            .DIN(N__12092),
            .DOUT(N__12091),
            .PACKAGEPIN(LMBEn));
    defparam LMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LMBEn_obuf_preio (
            .PADOEN(N__12093),
            .PADOUT(N__12092),
            .PADIN(N__12091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9413),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_11_iopad (
            .OE(N__12084),
            .DIN(N__12083),
            .DOUT(N__12082),
            .PACKAGEPIN(A[11]));
    defparam A_ibuf_11_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_11_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_11_preio (
            .PADOEN(N__12084),
            .PADOUT(N__12083),
            .PADIN(N__12082),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_11),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CUUBEn_obuf_iopad (
            .OE(N__12075),
            .DIN(N__12074),
            .DOUT(N__12073),
            .PACKAGEPIN(CUUBEn));
    defparam CUUBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CUUBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CUUBEn_obuf_preio (
            .PADOEN(N__12075),
            .PADOUT(N__12074),
            .PADIN(N__12073),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9551),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD TACKn_obuft_iopad (
            .OE(N__12066),
            .DIN(N__12065),
            .DOUT(N__12064),
            .PACKAGEPIN(TACKn));
    defparam TACKn_obuft_preio.NEG_TRIGGER=1'b0;
    defparam TACKn_obuft_preio.PIN_TYPE=6'b101001;
    PRE_IO TACKn_obuft_preio (
            .PADOEN(N__12066),
            .PADOUT(N__12065),
            .PADIN(N__12064),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__4461),
            .DIN0(),
            .DOUT0(N__5241),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_2_iopad (
            .OE(N__12057),
            .DIN(N__12056),
            .DOUT(N__12055),
            .PACKAGEPIN(CMA[2]));
    defparam CMA_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_2_preio (
            .PADOEN(N__12057),
            .PADOUT(N__12056),
            .PADIN(N__12055),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5330),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_4_iopad (
            .OE(N__12048),
            .DIN(N__12047),
            .DOUT(N__12046),
            .PACKAGEPIN(DRA[4]));
    defparam DRA_ibuf_4_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_4_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_4_preio (
            .PADOEN(N__12048),
            .PADOUT(N__12047),
            .PADIN(N__12046),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_14_iopad (
            .OE(N__12039),
            .DIN(N__12038),
            .DOUT(N__12037),
            .PACKAGEPIN(A[14]));
    defparam A_ibuf_14_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_14_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_14_preio (
            .PADOEN(N__12039),
            .PADOUT(N__12038),
            .PADIN(N__12037),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_14),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_8_iopad (
            .OE(N__12030),
            .DIN(N__12029),
            .DOUT(N__12028),
            .PACKAGEPIN(CMA[8]));
    defparam CMA_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_8_preio (
            .PADOEN(N__12030),
            .PADOUT(N__12029),
            .PADIN(N__12028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4652),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD AWEn_ibuf_iopad (
            .OE(N__12021),
            .DIN(N__12020),
            .DOUT(N__12019),
            .PACKAGEPIN(AWEn));
    defparam AWEn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam AWEn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO AWEn_ibuf_preio (
            .PADOEN(N__12021),
            .PADOUT(N__12020),
            .PADIN(N__12019),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(AWEn_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_1_iopad (
            .OE(N__12012),
            .DIN(N__12011),
            .DOUT(N__12010),
            .PACKAGEPIN(DRA[1]));
    defparam DRA_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_1_preio (
            .PADOEN(N__12012),
            .PADOUT(N__12011),
            .PADIN(N__12010),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DA_obuf_1_iopad (
            .OE(N__12003),
            .DIN(N__12002),
            .DOUT(N__12001),
            .PACKAGEPIN(DA[1]));
    defparam DA_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam DA_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO DA_obuf_1_preio (
            .PADOEN(N__12003),
            .PADOUT(N__12002),
            .PADIN(N__12001),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4730),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_17_iopad (
            .OE(N__11994),
            .DIN(N__11993),
            .DOUT(N__11992),
            .PACKAGEPIN(A[17]));
    defparam A_ibuf_17_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_17_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_17_preio (
            .PADOEN(N__11994),
            .PADOUT(N__11993),
            .PADIN(N__11992),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_17),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_1_iopad (
            .OE(N__11985),
            .DIN(N__11984),
            .DOUT(N__11983),
            .PACKAGEPIN(A[1]));
    defparam A_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_1_preio (
            .PADOEN(N__11985),
            .PADOUT(N__11984),
            .PADIN(N__11983),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_5_iopad (
            .OE(N__11976),
            .DIN(N__11975),
            .DOUT(N__11974),
            .PACKAGEPIN(CMA[5]));
    defparam CMA_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_5_preio (
            .PADOEN(N__11976),
            .PADOUT(N__11975),
            .PADIN(N__11974),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4529),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UDSn_obuf_iopad (
            .OE(N__11967),
            .DIN(N__11966),
            .DOUT(N__11965),
            .PACKAGEPIN(UDSn));
    defparam UDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UDSn_obuf_preio (
            .PADOEN(N__11967),
            .PADOUT(N__11966),
            .PADIN(N__11965),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8672),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD UMBEn_obuf_iopad (
            .OE(N__11958),
            .DIN(N__11957),
            .DOUT(N__11956),
            .PACKAGEPIN(UMBEn));
    defparam UMBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam UMBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO UMBEn_obuf_preio (
            .PADOEN(N__11958),
            .PADOUT(N__11957),
            .PADIN(N__11956),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11288),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK_EN_obuf_iopad (
            .OE(N__11949),
            .DIN(N__11948),
            .DOUT(N__11947),
            .PACKAGEPIN(CLK_EN));
    defparam CLK_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK_EN_obuf_preio (
            .PADOEN(N__11949),
            .PADOUT(N__11948),
            .PADIN(N__11947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5717),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_2_iopad (
            .OE(N__11940),
            .DIN(N__11939),
            .DOUT(N__11938),
            .PACKAGEPIN(DRA[2]));
    defparam DRA_ibuf_2_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_2_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_2_preio (
            .PADOEN(N__11940),
            .PADOUT(N__11939),
            .PADIN(N__11938),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_6_iopad (
            .OE(N__11931),
            .DIN(N__11930),
            .DOUT(N__11929),
            .PACKAGEPIN(A[6]));
    defparam A_ibuf_6_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_6_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_6_preio (
            .PADOEN(N__11931),
            .PADOUT(N__11930),
            .PADIN(N__11929),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_6_iopad (
            .OE(N__11922),
            .DIN(N__11921),
            .DOUT(N__11920),
            .PACKAGEPIN(CMA[6]));
    defparam CMA_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_6_preio (
            .PADOEN(N__11922),
            .PADOUT(N__11921),
            .PADIN(N__11920),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8459),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_8_iopad (
            .OE(N__11913),
            .DIN(N__11912),
            .DOUT(N__11911),
            .PACKAGEPIN(DRA[8]));
    defparam DRA_ibuf_8_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_8_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_8_preio (
            .PADOEN(N__11913),
            .PADOUT(N__11912),
            .PADIN(N__11911),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_10_iopad (
            .OE(N__11904),
            .DIN(N__11903),
            .DOUT(N__11902),
            .PACKAGEPIN(A[10]));
    defparam A_ibuf_10_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_10_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_10_preio (
            .PADOEN(N__11904),
            .PADOUT(N__11903),
            .PADIN(N__11902),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_10),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LATCH_CLK_obuf_iopad (
            .OE(N__11895),
            .DIN(N__11894),
            .DOUT(N__11893),
            .PACKAGEPIN(LATCH_CLK));
    defparam LATCH_CLK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LATCH_CLK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LATCH_CLK_obuf_preio (
            .PADOEN(N__11895),
            .PADOUT(N__11894),
            .PADIN(N__11893),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5048),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LDSn_obuf_iopad (
            .OE(N__11886),
            .DIN(N__11885),
            .DOUT(N__11884),
            .PACKAGEPIN(LDSn));
    defparam LDSn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LDSn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LDSn_obuf_preio (
            .PADOEN(N__11886),
            .PADOUT(N__11885),
            .PADIN(N__11884),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8174),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40B_OUT_obuf_iopad (
            .OE(N__11877),
            .DIN(N__11876),
            .DOUT(N__11875),
            .PACKAGEPIN(CLK40B_OUT));
    defparam CLK40B_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40B_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40B_OUT_obuf_preio (
            .PADOEN(N__11877),
            .PADOUT(N__11876),
            .PADIN(N__11875),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9482),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SIZ_ibuf_1_iopad (
            .OE(N__11868),
            .DIN(N__11867),
            .DOUT(N__11866),
            .PACKAGEPIN(SIZ[1]));
    defparam SIZ_ibuf_1_preio.NEG_TRIGGER=1'b0;
    defparam SIZ_ibuf_1_preio.PIN_TYPE=6'b000001;
    PRE_IO SIZ_ibuf_1_preio (
            .PADOEN(N__11868),
            .PADOUT(N__11867),
            .PADIN(N__11866),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SIZ_c_1),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40D_OUT_obuf_iopad (
            .OE(N__11859),
            .DIN(N__11858),
            .DOUT(N__11857),
            .PACKAGEPIN(CLK40D_OUT));
    defparam CLK40D_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40D_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40D_OUT_obuf_preio (
            .PADOEN(N__11859),
            .PADOUT(N__11858),
            .PADIN(N__11857),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9471),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLKRAM_obuf_iopad (
            .OE(N__11850),
            .DIN(N__11849),
            .DOUT(N__11848),
            .PACKAGEPIN(CLKRAM));
    defparam CLKRAM_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLKRAM_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLKRAM_obuf_preio (
            .PADOEN(N__11850),
            .PADOUT(N__11849),
            .PADIN(N__11848),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4430),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_3_iopad (
            .OE(N__11841),
            .DIN(N__11840),
            .DOUT(N__11839),
            .PACKAGEPIN(CMA[3]));
    defparam CMA_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_3_preio (
            .PADOEN(N__11841),
            .PADOUT(N__11840),
            .PADIN(N__11839),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8618),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_20_iopad (
            .OE(N__11832),
            .DIN(N__11831),
            .DOUT(N__11830),
            .PACKAGEPIN(A[20]));
    defparam A_ibuf_20_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_20_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_20_preio (
            .PADOEN(N__11832),
            .PADOUT(N__11831),
            .PADIN(N__11830),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_20),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD C3_ibuf_iopad (
            .OE(N__11823),
            .DIN(N__11822),
            .DOUT(N__11821),
            .PACKAGEPIN(C3));
    defparam C3_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam C3_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO C3_ibuf_preio (
            .PADOEN(N__11823),
            .PADOUT(N__11822),
            .PADIN(N__11821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(C3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRA_ibuf_5_iopad (
            .OE(N__11814),
            .DIN(N__11813),
            .DOUT(N__11812),
            .PACKAGEPIN(DRA[5]));
    defparam DRA_ibuf_5_preio.NEG_TRIGGER=1'b0;
    defparam DRA_ibuf_5_preio.PIN_TYPE=6'b000001;
    PRE_IO DRA_ibuf_5_preio (
            .PADOEN(N__11814),
            .PADOUT(N__11813),
            .PADIN(N__11812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DRA_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD A_ibuf_13_iopad (
            .OE(N__11805),
            .DIN(N__11804),
            .DOUT(N__11803),
            .PACKAGEPIN(A[13]));
    defparam A_ibuf_13_preio.NEG_TRIGGER=1'b0;
    defparam A_ibuf_13_preio.PIN_TYPE=6'b000001;
    PRE_IO A_ibuf_13_preio (
            .PADOEN(N__11805),
            .PADOUT(N__11804),
            .PADIN(N__11803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(A_c_13),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLK40C_OUT_obuf_iopad (
            .OE(N__11796),
            .DIN(N__11795),
            .DOUT(N__11794),
            .PACKAGEPIN(CLK40C_OUT));
    defparam CLK40C_OUT_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLK40C_OUT_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLK40C_OUT_obuf_preio (
            .PADOEN(N__11796),
            .PADOUT(N__11795),
            .PADIN(N__11794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DRDENn_obuf_iopad (
            .OE(N__11787),
            .DIN(N__11786),
            .DOUT(N__11785),
            .PACKAGEPIN(DRDENn));
    defparam DRDENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DRDENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DRDENn_obuf_preio (
            .PADOEN(N__11787),
            .PADOUT(N__11786),
            .PADIN(N__11785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9917),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CLLBEn_obuf_iopad (
            .OE(N__11778),
            .DIN(N__11777),
            .DOUT(N__11776),
            .PACKAGEPIN(CLLBEn));
    defparam CLLBEn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam CLLBEn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO CLLBEn_obuf_preio (
            .PADOEN(N__11778),
            .PADOUT(N__11777),
            .PADIN(N__11776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8393),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD CMA_obuf_9_iopad (
            .OE(N__11769),
            .DIN(N__11768),
            .DOUT(N__11767),
            .PACKAGEPIN(CMA[9]));
    defparam CMA_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam CMA_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO CMA_obuf_9_preio (
            .PADOEN(N__11769),
            .PADOUT(N__11768),
            .PADIN(N__11767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2838 (
            .O(N__11750),
            .I(N__11745));
    InMux I__2837 (
            .O(N__11749),
            .I(N__11738));
    InMux I__2836 (
            .O(N__11748),
            .I(N__11738));
    LocalMux I__2835 (
            .O(N__11745),
            .I(N__11735));
    InMux I__2834 (
            .O(N__11744),
            .I(N__11732));
    CascadeMux I__2833 (
            .O(N__11743),
            .I(N__11728));
    LocalMux I__2832 (
            .O(N__11738),
            .I(N__11725));
    Sp12to4 I__2831 (
            .O(N__11735),
            .I(N__11722));
    LocalMux I__2830 (
            .O(N__11732),
            .I(N__11719));
    InMux I__2829 (
            .O(N__11731),
            .I(N__11716));
    InMux I__2828 (
            .O(N__11728),
            .I(N__11713));
    Span12Mux_h I__2827 (
            .O(N__11725),
            .I(N__11710));
    Span12Mux_v I__2826 (
            .O(N__11722),
            .I(N__11707));
    Span12Mux_h I__2825 (
            .O(N__11719),
            .I(N__11700));
    LocalMux I__2824 (
            .O(N__11716),
            .I(N__11700));
    LocalMux I__2823 (
            .O(N__11713),
            .I(N__11700));
    Span12Mux_v I__2822 (
            .O(N__11710),
            .I(N__11697));
    Span12Mux_h I__2821 (
            .O(N__11707),
            .I(N__11692));
    Span12Mux_v I__2820 (
            .O(N__11700),
            .I(N__11692));
    Odrv12 I__2819 (
            .O(N__11697),
            .I(CASLn_c));
    Odrv12 I__2818 (
            .O(N__11692),
            .I(CASLn_c));
    InMux I__2817 (
            .O(N__11687),
            .I(N__11684));
    LocalMux I__2816 (
            .O(N__11684),
            .I(N__11681));
    Span4Mux_v I__2815 (
            .O(N__11681),
            .I(N__11678));
    Sp12to4 I__2814 (
            .O(N__11678),
            .I(N__11674));
    InMux I__2813 (
            .O(N__11677),
            .I(N__11671));
    Span12Mux_h I__2812 (
            .O(N__11674),
            .I(N__11665));
    LocalMux I__2811 (
            .O(N__11671),
            .I(N__11665));
    CascadeMux I__2810 (
            .O(N__11670),
            .I(N__11662));
    Span12Mux_s11_v I__2809 (
            .O(N__11665),
            .I(N__11659));
    InMux I__2808 (
            .O(N__11662),
            .I(N__11656));
    Odrv12 I__2807 (
            .O(N__11659),
            .I(DMA_WRITE_CYCLE));
    LocalMux I__2806 (
            .O(N__11656),
            .I(DMA_WRITE_CYCLE));
    IoInMux I__2805 (
            .O(N__11651),
            .I(N__11648));
    LocalMux I__2804 (
            .O(N__11648),
            .I(N__11645));
    IoSpan4Mux I__2803 (
            .O(N__11645),
            .I(N__11642));
    Span4Mux_s3_v I__2802 (
            .O(N__11642),
            .I(N__11639));
    Span4Mux_v I__2801 (
            .O(N__11639),
            .I(N__11636));
    Odrv4 I__2800 (
            .O(N__11636),
            .I(N_357));
    IoInMux I__2799 (
            .O(N__11633),
            .I(N__11630));
    LocalMux I__2798 (
            .O(N__11630),
            .I(N__11627));
    Span4Mux_s3_v I__2797 (
            .O(N__11627),
            .I(N__11624));
    Odrv4 I__2796 (
            .O(N__11624),
            .I(N_373_i));
    InMux I__2795 (
            .O(N__11621),
            .I(N__11615));
    InMux I__2794 (
            .O(N__11620),
            .I(N__11615));
    LocalMux I__2793 (
            .O(N__11615),
            .I(N__11606));
    InMux I__2792 (
            .O(N__11614),
            .I(N__11599));
    InMux I__2791 (
            .O(N__11613),
            .I(N__11599));
    InMux I__2790 (
            .O(N__11612),
            .I(N__11599));
    InMux I__2789 (
            .O(N__11611),
            .I(N__11596));
    InMux I__2788 (
            .O(N__11610),
            .I(N__11591));
    InMux I__2787 (
            .O(N__11609),
            .I(N__11591));
    Span4Mux_v I__2786 (
            .O(N__11606),
            .I(N__11588));
    LocalMux I__2785 (
            .O(N__11599),
            .I(N__11585));
    LocalMux I__2784 (
            .O(N__11596),
            .I(N__11582));
    LocalMux I__2783 (
            .O(N__11591),
            .I(N__11579));
    Span4Mux_v I__2782 (
            .O(N__11588),
            .I(N__11574));
    Span4Mux_v I__2781 (
            .O(N__11585),
            .I(N__11574));
    Span4Mux_v I__2780 (
            .O(N__11582),
            .I(N__11571));
    Span12Mux_v I__2779 (
            .O(N__11579),
            .I(N__11568));
    Sp12to4 I__2778 (
            .O(N__11574),
            .I(N__11563));
    Sp12to4 I__2777 (
            .O(N__11571),
            .I(N__11563));
    Span12Mux_h I__2776 (
            .O(N__11568),
            .I(N__11560));
    Span12Mux_h I__2775 (
            .O(N__11563),
            .I(N__11557));
    Odrv12 I__2774 (
            .O(N__11560),
            .I(A_c_1));
    Odrv12 I__2773 (
            .O(N__11557),
            .I(A_c_1));
    InMux I__2772 (
            .O(N__11552),
            .I(N__11540));
    InMux I__2771 (
            .O(N__11551),
            .I(N__11540));
    InMux I__2770 (
            .O(N__11550),
            .I(N__11540));
    InMux I__2769 (
            .O(N__11549),
            .I(N__11535));
    InMux I__2768 (
            .O(N__11548),
            .I(N__11535));
    InMux I__2767 (
            .O(N__11547),
            .I(N__11531));
    LocalMux I__2766 (
            .O(N__11540),
            .I(N__11527));
    LocalMux I__2765 (
            .O(N__11535),
            .I(N__11524));
    InMux I__2764 (
            .O(N__11534),
            .I(N__11521));
    LocalMux I__2763 (
            .O(N__11531),
            .I(N__11518));
    InMux I__2762 (
            .O(N__11530),
            .I(N__11515));
    Span4Mux_v I__2761 (
            .O(N__11527),
            .I(N__11510));
    Span4Mux_v I__2760 (
            .O(N__11524),
            .I(N__11510));
    LocalMux I__2759 (
            .O(N__11521),
            .I(N__11507));
    Span4Mux_v I__2758 (
            .O(N__11518),
            .I(N__11503));
    LocalMux I__2757 (
            .O(N__11515),
            .I(N__11500));
    Span4Mux_h I__2756 (
            .O(N__11510),
            .I(N__11495));
    Span4Mux_v I__2755 (
            .O(N__11507),
            .I(N__11495));
    InMux I__2754 (
            .O(N__11506),
            .I(N__11492));
    Sp12to4 I__2753 (
            .O(N__11503),
            .I(N__11487));
    Span12Mux_v I__2752 (
            .O(N__11500),
            .I(N__11487));
    Sp12to4 I__2751 (
            .O(N__11495),
            .I(N__11482));
    LocalMux I__2750 (
            .O(N__11492),
            .I(N__11482));
    Span12Mux_h I__2749 (
            .O(N__11487),
            .I(N__11479));
    Span12Mux_h I__2748 (
            .O(N__11482),
            .I(N__11476));
    Odrv12 I__2747 (
            .O(N__11479),
            .I(A_c_0));
    Odrv12 I__2746 (
            .O(N__11476),
            .I(A_c_0));
    InMux I__2745 (
            .O(N__11471),
            .I(N__11467));
    InMux I__2744 (
            .O(N__11470),
            .I(N__11459));
    LocalMux I__2743 (
            .O(N__11467),
            .I(N__11456));
    InMux I__2742 (
            .O(N__11466),
            .I(N__11453));
    InMux I__2741 (
            .O(N__11465),
            .I(N__11450));
    CascadeMux I__2740 (
            .O(N__11464),
            .I(N__11447));
    CascadeMux I__2739 (
            .O(N__11463),
            .I(N__11444));
    CascadeMux I__2738 (
            .O(N__11462),
            .I(N__11441));
    LocalMux I__2737 (
            .O(N__11459),
            .I(N__11437));
    Span4Mux_v I__2736 (
            .O(N__11456),
            .I(N__11432));
    LocalMux I__2735 (
            .O(N__11453),
            .I(N__11432));
    LocalMux I__2734 (
            .O(N__11450),
            .I(N__11429));
    InMux I__2733 (
            .O(N__11447),
            .I(N__11422));
    InMux I__2732 (
            .O(N__11444),
            .I(N__11422));
    InMux I__2731 (
            .O(N__11441),
            .I(N__11422));
    InMux I__2730 (
            .O(N__11440),
            .I(N__11419));
    Span4Mux_v I__2729 (
            .O(N__11437),
            .I(N__11416));
    Span4Mux_h I__2728 (
            .O(N__11432),
            .I(N__11411));
    Span4Mux_v I__2727 (
            .O(N__11429),
            .I(N__11411));
    LocalMux I__2726 (
            .O(N__11422),
            .I(N__11406));
    LocalMux I__2725 (
            .O(N__11419),
            .I(N__11406));
    Span4Mux_v I__2724 (
            .O(N__11416),
            .I(N__11403));
    Span4Mux_v I__2723 (
            .O(N__11411),
            .I(N__11398));
    Span4Mux_h I__2722 (
            .O(N__11406),
            .I(N__11398));
    Span4Mux_v I__2721 (
            .O(N__11403),
            .I(N__11395));
    Span4Mux_v I__2720 (
            .O(N__11398),
            .I(N__11392));
    Sp12to4 I__2719 (
            .O(N__11395),
            .I(N__11387));
    Sp12to4 I__2718 (
            .O(N__11392),
            .I(N__11387));
    Span12Mux_h I__2717 (
            .O(N__11387),
            .I(N__11384));
    Odrv12 I__2716 (
            .O(N__11384),
            .I(SIZ_c_0));
    CascadeMux I__2715 (
            .O(N__11381),
            .I(N__11376));
    InMux I__2714 (
            .O(N__11380),
            .I(N__11372));
    InMux I__2713 (
            .O(N__11379),
            .I(N__11369));
    InMux I__2712 (
            .O(N__11376),
            .I(N__11366));
    InMux I__2711 (
            .O(N__11375),
            .I(N__11363));
    LocalMux I__2710 (
            .O(N__11372),
            .I(N__11357));
    LocalMux I__2709 (
            .O(N__11369),
            .I(N__11357));
    LocalMux I__2708 (
            .O(N__11366),
            .I(N__11354));
    LocalMux I__2707 (
            .O(N__11363),
            .I(N__11351));
    CascadeMux I__2706 (
            .O(N__11362),
            .I(N__11345));
    Span4Mux_v I__2705 (
            .O(N__11357),
            .I(N__11342));
    Span4Mux_h I__2704 (
            .O(N__11354),
            .I(N__11337));
    Span4Mux_v I__2703 (
            .O(N__11351),
            .I(N__11337));
    InMux I__2702 (
            .O(N__11350),
            .I(N__11329));
    InMux I__2701 (
            .O(N__11349),
            .I(N__11329));
    InMux I__2700 (
            .O(N__11348),
            .I(N__11329));
    InMux I__2699 (
            .O(N__11345),
            .I(N__11326));
    Span4Mux_v I__2698 (
            .O(N__11342),
            .I(N__11323));
    Span4Mux_v I__2697 (
            .O(N__11337),
            .I(N__11320));
    InMux I__2696 (
            .O(N__11336),
            .I(N__11317));
    LocalMux I__2695 (
            .O(N__11329),
            .I(N__11312));
    LocalMux I__2694 (
            .O(N__11326),
            .I(N__11312));
    Span4Mux_v I__2693 (
            .O(N__11323),
            .I(N__11309));
    Span4Mux_v I__2692 (
            .O(N__11320),
            .I(N__11306));
    LocalMux I__2691 (
            .O(N__11317),
            .I(N__11301));
    Sp12to4 I__2690 (
            .O(N__11312),
            .I(N__11301));
    Sp12to4 I__2689 (
            .O(N__11309),
            .I(N__11294));
    Sp12to4 I__2688 (
            .O(N__11306),
            .I(N__11294));
    Span12Mux_v I__2687 (
            .O(N__11301),
            .I(N__11294));
    Span12Mux_h I__2686 (
            .O(N__11294),
            .I(N__11291));
    Odrv12 I__2685 (
            .O(N__11291),
            .I(SIZ_c_1));
    IoInMux I__2684 (
            .O(N__11288),
            .I(N__11285));
    LocalMux I__2683 (
            .O(N__11285),
            .I(N__11282));
    Span4Mux_s2_v I__2682 (
            .O(N__11282),
            .I(N__11279));
    Span4Mux_h I__2681 (
            .O(N__11279),
            .I(N__11276));
    Span4Mux_v I__2680 (
            .O(N__11276),
            .I(N__11273));
    Odrv4 I__2679 (
            .O(N__11273),
            .I(UMBEn_c));
    InMux I__2678 (
            .O(N__11270),
            .I(N__11267));
    LocalMux I__2677 (
            .O(N__11267),
            .I(N__11264));
    Odrv12 I__2676 (
            .O(N__11264),
            .I(\U712_CHIP_RAM.CMA_5_i_0_9 ));
    InMux I__2675 (
            .O(N__11261),
            .I(N__11258));
    LocalMux I__2674 (
            .O(N__11258),
            .I(N__11255));
    Sp12to4 I__2673 (
            .O(N__11255),
            .I(N__11252));
    Span12Mux_v I__2672 (
            .O(N__11252),
            .I(N__11249));
    Span12Mux_h I__2671 (
            .O(N__11249),
            .I(N__11246));
    Odrv12 I__2670 (
            .O(N__11246),
            .I(A_c_19));
    IoInMux I__2669 (
            .O(N__11243),
            .I(N__11240));
    LocalMux I__2668 (
            .O(N__11240),
            .I(N__11237));
    IoSpan4Mux I__2667 (
            .O(N__11237),
            .I(N__11234));
    IoSpan4Mux I__2666 (
            .O(N__11234),
            .I(N__11231));
    Span4Mux_s2_h I__2665 (
            .O(N__11231),
            .I(N__11228));
    Sp12to4 I__2664 (
            .O(N__11228),
            .I(N__11225));
    Odrv12 I__2663 (
            .O(N__11225),
            .I(CMA_c_9));
    CEMux I__2662 (
            .O(N__11222),
            .I(N__11219));
    LocalMux I__2661 (
            .O(N__11219),
            .I(N__11214));
    CEMux I__2660 (
            .O(N__11218),
            .I(N__11211));
    CEMux I__2659 (
            .O(N__11217),
            .I(N__11208));
    Span4Mux_v I__2658 (
            .O(N__11214),
            .I(N__11202));
    LocalMux I__2657 (
            .O(N__11211),
            .I(N__11202));
    LocalMux I__2656 (
            .O(N__11208),
            .I(N__11199));
    CEMux I__2655 (
            .O(N__11207),
            .I(N__11196));
    Sp12to4 I__2654 (
            .O(N__11202),
            .I(N__11192));
    Span4Mux_h I__2653 (
            .O(N__11199),
            .I(N__11187));
    LocalMux I__2652 (
            .O(N__11196),
            .I(N__11187));
    CEMux I__2651 (
            .O(N__11195),
            .I(N__11184));
    Span12Mux_h I__2650 (
            .O(N__11192),
            .I(N__11179));
    Sp12to4 I__2649 (
            .O(N__11187),
            .I(N__11179));
    LocalMux I__2648 (
            .O(N__11184),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    Odrv12 I__2647 (
            .O(N__11179),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_0 ));
    CascadeMux I__2646 (
            .O(N__11174),
            .I(N__11169));
    InMux I__2645 (
            .O(N__11173),
            .I(N__11165));
    InMux I__2644 (
            .O(N__11172),
            .I(N__11160));
    InMux I__2643 (
            .O(N__11169),
            .I(N__11157));
    InMux I__2642 (
            .O(N__11168),
            .I(N__11154));
    LocalMux I__2641 (
            .O(N__11165),
            .I(N__11150));
    InMux I__2640 (
            .O(N__11164),
            .I(N__11147));
    InMux I__2639 (
            .O(N__11163),
            .I(N__11144));
    LocalMux I__2638 (
            .O(N__11160),
            .I(N__11141));
    LocalMux I__2637 (
            .O(N__11157),
            .I(N__11138));
    LocalMux I__2636 (
            .O(N__11154),
            .I(N__11135));
    InMux I__2635 (
            .O(N__11153),
            .I(N__11132));
    Span4Mux_h I__2634 (
            .O(N__11150),
            .I(N__11126));
    LocalMux I__2633 (
            .O(N__11147),
            .I(N__11126));
    LocalMux I__2632 (
            .O(N__11144),
            .I(N__11123));
    Span4Mux_v I__2631 (
            .O(N__11141),
            .I(N__11118));
    Span4Mux_v I__2630 (
            .O(N__11138),
            .I(N__11118));
    Span4Mux_h I__2629 (
            .O(N__11135),
            .I(N__11113));
    LocalMux I__2628 (
            .O(N__11132),
            .I(N__11113));
    InMux I__2627 (
            .O(N__11131),
            .I(N__11110));
    Odrv4 I__2626 (
            .O(N__11126),
            .I(DMA_CYCLEm));
    Odrv4 I__2625 (
            .O(N__11123),
            .I(DMA_CYCLEm));
    Odrv4 I__2624 (
            .O(N__11118),
            .I(DMA_CYCLEm));
    Odrv4 I__2623 (
            .O(N__11113),
            .I(DMA_CYCLEm));
    LocalMux I__2622 (
            .O(N__11110),
            .I(DMA_CYCLEm));
    InMux I__2621 (
            .O(N__11099),
            .I(N__11096));
    LocalMux I__2620 (
            .O(N__11096),
            .I(\U712_BYTE_ENABLE.N_411 ));
    IoInMux I__2619 (
            .O(N__11093),
            .I(N__11090));
    LocalMux I__2618 (
            .O(N__11090),
            .I(N__11085));
    InMux I__2617 (
            .O(N__11089),
            .I(N__11082));
    InMux I__2616 (
            .O(N__11088),
            .I(N__11079));
    Span4Mux_s2_v I__2615 (
            .O(N__11085),
            .I(N__11075));
    LocalMux I__2614 (
            .O(N__11082),
            .I(N__11072));
    LocalMux I__2613 (
            .O(N__11079),
            .I(N__11069));
    InMux I__2612 (
            .O(N__11078),
            .I(N__11066));
    Span4Mux_v I__2611 (
            .O(N__11075),
            .I(N__11063));
    Span4Mux_v I__2610 (
            .O(N__11072),
            .I(N__11059));
    Span4Mux_v I__2609 (
            .O(N__11069),
            .I(N__11056));
    LocalMux I__2608 (
            .O(N__11066),
            .I(N__11053));
    Sp12to4 I__2607 (
            .O(N__11063),
            .I(N__11050));
    InMux I__2606 (
            .O(N__11062),
            .I(N__11047));
    Span4Mux_v I__2605 (
            .O(N__11059),
            .I(N__11043));
    Span4Mux_h I__2604 (
            .O(N__11056),
            .I(N__11038));
    Span4Mux_v I__2603 (
            .O(N__11053),
            .I(N__11038));
    Span12Mux_h I__2602 (
            .O(N__11050),
            .I(N__11033));
    LocalMux I__2601 (
            .O(N__11047),
            .I(N__11033));
    InMux I__2600 (
            .O(N__11046),
            .I(N__11030));
    Odrv4 I__2599 (
            .O(N__11043),
            .I(DBENn_c));
    Odrv4 I__2598 (
            .O(N__11038),
            .I(DBENn_c));
    Odrv12 I__2597 (
            .O(N__11033),
            .I(DBENn_c));
    LocalMux I__2596 (
            .O(N__11030),
            .I(DBENn_c));
    IoInMux I__2595 (
            .O(N__11021),
            .I(N__11018));
    LocalMux I__2594 (
            .O(N__11018),
            .I(N__11015));
    Span4Mux_s1_h I__2593 (
            .O(N__11015),
            .I(N__11012));
    Sp12to4 I__2592 (
            .O(N__11012),
            .I(N__11009));
    Span12Mux_v I__2591 (
            .O(N__11009),
            .I(N__11006));
    Span12Mux_h I__2590 (
            .O(N__11006),
            .I(N__11003));
    Odrv12 I__2589 (
            .O(N__11003),
            .I(N_150_i));
    CascadeMux I__2588 (
            .O(N__11000),
            .I(N__10991));
    CascadeMux I__2587 (
            .O(N__10999),
            .I(N__10987));
    CascadeMux I__2586 (
            .O(N__10998),
            .I(N__10984));
    CascadeMux I__2585 (
            .O(N__10997),
            .I(N__10975));
    InMux I__2584 (
            .O(N__10996),
            .I(N__10972));
    InMux I__2583 (
            .O(N__10995),
            .I(N__10969));
    InMux I__2582 (
            .O(N__10994),
            .I(N__10954));
    InMux I__2581 (
            .O(N__10991),
            .I(N__10954));
    InMux I__2580 (
            .O(N__10990),
            .I(N__10954));
    InMux I__2579 (
            .O(N__10987),
            .I(N__10954));
    InMux I__2578 (
            .O(N__10984),
            .I(N__10954));
    InMux I__2577 (
            .O(N__10983),
            .I(N__10954));
    InMux I__2576 (
            .O(N__10982),
            .I(N__10954));
    InMux I__2575 (
            .O(N__10981),
            .I(N__10949));
    InMux I__2574 (
            .O(N__10980),
            .I(N__10949));
    InMux I__2573 (
            .O(N__10979),
            .I(N__10946));
    InMux I__2572 (
            .O(N__10978),
            .I(N__10942));
    InMux I__2571 (
            .O(N__10975),
            .I(N__10939));
    LocalMux I__2570 (
            .O(N__10972),
            .I(N__10924));
    LocalMux I__2569 (
            .O(N__10969),
            .I(N__10924));
    LocalMux I__2568 (
            .O(N__10954),
            .I(N__10924));
    LocalMux I__2567 (
            .O(N__10949),
            .I(N__10924));
    LocalMux I__2566 (
            .O(N__10946),
            .I(N__10921));
    InMux I__2565 (
            .O(N__10945),
            .I(N__10918));
    LocalMux I__2564 (
            .O(N__10942),
            .I(N__10915));
    LocalMux I__2563 (
            .O(N__10939),
            .I(N__10912));
    InMux I__2562 (
            .O(N__10938),
            .I(N__10905));
    InMux I__2561 (
            .O(N__10937),
            .I(N__10905));
    InMux I__2560 (
            .O(N__10936),
            .I(N__10905));
    InMux I__2559 (
            .O(N__10935),
            .I(N__10902));
    InMux I__2558 (
            .O(N__10934),
            .I(N__10899));
    InMux I__2557 (
            .O(N__10933),
            .I(N__10896));
    Span4Mux_v I__2556 (
            .O(N__10924),
            .I(N__10889));
    Span4Mux_h I__2555 (
            .O(N__10921),
            .I(N__10889));
    LocalMux I__2554 (
            .O(N__10918),
            .I(N__10889));
    Span4Mux_v I__2553 (
            .O(N__10915),
            .I(N__10886));
    Span12Mux_h I__2552 (
            .O(N__10912),
            .I(N__10879));
    LocalMux I__2551 (
            .O(N__10905),
            .I(N__10879));
    LocalMux I__2550 (
            .O(N__10902),
            .I(N__10879));
    LocalMux I__2549 (
            .O(N__10899),
            .I(N__10872));
    LocalMux I__2548 (
            .O(N__10896),
            .I(N__10872));
    Sp12to4 I__2547 (
            .O(N__10889),
            .I(N__10872));
    Sp12to4 I__2546 (
            .O(N__10886),
            .I(N__10869));
    Span12Mux_h I__2545 (
            .O(N__10879),
            .I(N__10866));
    Span12Mux_v I__2544 (
            .O(N__10872),
            .I(N__10863));
    Span12Mux_h I__2543 (
            .O(N__10869),
            .I(N__10860));
    Span12Mux_v I__2542 (
            .O(N__10866),
            .I(N__10855));
    Span12Mux_h I__2541 (
            .O(N__10863),
            .I(N__10855));
    Span12Mux_v I__2540 (
            .O(N__10860),
            .I(N__10852));
    Odrv12 I__2539 (
            .O(N__10855),
            .I(AGNUS_REV_c));
    Odrv12 I__2538 (
            .O(N__10852),
            .I(AGNUS_REV_c));
    CascadeMux I__2537 (
            .O(N__10847),
            .I(N__10842));
    InMux I__2536 (
            .O(N__10846),
            .I(N__10839));
    InMux I__2535 (
            .O(N__10845),
            .I(N__10836));
    InMux I__2534 (
            .O(N__10842),
            .I(N__10833));
    LocalMux I__2533 (
            .O(N__10839),
            .I(N__10829));
    LocalMux I__2532 (
            .O(N__10836),
            .I(N__10824));
    LocalMux I__2531 (
            .O(N__10833),
            .I(N__10824));
    InMux I__2530 (
            .O(N__10832),
            .I(N__10821));
    Span4Mux_h I__2529 (
            .O(N__10829),
            .I(N__10814));
    Span4Mux_v I__2528 (
            .O(N__10824),
            .I(N__10814));
    LocalMux I__2527 (
            .O(N__10821),
            .I(N__10814));
    Span4Mux_h I__2526 (
            .O(N__10814),
            .I(N__10811));
    Span4Mux_v I__2525 (
            .O(N__10811),
            .I(N__10808));
    Sp12to4 I__2524 (
            .O(N__10808),
            .I(N__10805));
    Span12Mux_v I__2523 (
            .O(N__10805),
            .I(N__10802));
    Odrv12 I__2522 (
            .O(N__10802),
            .I(DRA_c_9));
    InMux I__2521 (
            .O(N__10799),
            .I(N__10796));
    LocalMux I__2520 (
            .O(N__10796),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ));
    ClkMux I__2519 (
            .O(N__10793),
            .I(N__10775));
    ClkMux I__2518 (
            .O(N__10792),
            .I(N__10775));
    ClkMux I__2517 (
            .O(N__10791),
            .I(N__10775));
    ClkMux I__2516 (
            .O(N__10790),
            .I(N__10775));
    ClkMux I__2515 (
            .O(N__10789),
            .I(N__10775));
    ClkMux I__2514 (
            .O(N__10788),
            .I(N__10775));
    GlobalMux I__2513 (
            .O(N__10775),
            .I(N__10772));
    gio2CtrlBuf I__2512 (
            .O(N__10772),
            .I(C3_c_g));
    CEMux I__2511 (
            .O(N__10769),
            .I(N__10742));
    CEMux I__2510 (
            .O(N__10768),
            .I(N__10742));
    CEMux I__2509 (
            .O(N__10767),
            .I(N__10742));
    CEMux I__2508 (
            .O(N__10766),
            .I(N__10742));
    CEMux I__2507 (
            .O(N__10765),
            .I(N__10742));
    CEMux I__2506 (
            .O(N__10764),
            .I(N__10742));
    CEMux I__2505 (
            .O(N__10763),
            .I(N__10742));
    CEMux I__2504 (
            .O(N__10762),
            .I(N__10742));
    CEMux I__2503 (
            .O(N__10761),
            .I(N__10742));
    GlobalMux I__2502 (
            .O(N__10742),
            .I(N__10739));
    gio2CtrlBuf I__2501 (
            .O(N__10739),
            .I(DBRn_c_i_0_g));
    InMux I__2500 (
            .O(N__10736),
            .I(N__10726));
    InMux I__2499 (
            .O(N__10735),
            .I(N__10719));
    InMux I__2498 (
            .O(N__10734),
            .I(N__10719));
    InMux I__2497 (
            .O(N__10733),
            .I(N__10719));
    InMux I__2496 (
            .O(N__10732),
            .I(N__10716));
    InMux I__2495 (
            .O(N__10731),
            .I(N__10711));
    InMux I__2494 (
            .O(N__10730),
            .I(N__10711));
    InMux I__2493 (
            .O(N__10729),
            .I(N__10708));
    LocalMux I__2492 (
            .O(N__10726),
            .I(N__10704));
    LocalMux I__2491 (
            .O(N__10719),
            .I(N__10691));
    LocalMux I__2490 (
            .O(N__10716),
            .I(N__10683));
    LocalMux I__2489 (
            .O(N__10711),
            .I(N__10676));
    LocalMux I__2488 (
            .O(N__10708),
            .I(N__10658));
    SRMux I__2487 (
            .O(N__10707),
            .I(N__10574));
    Glb2LocalMux I__2486 (
            .O(N__10704),
            .I(N__10574));
    SRMux I__2485 (
            .O(N__10703),
            .I(N__10574));
    SRMux I__2484 (
            .O(N__10702),
            .I(N__10574));
    SRMux I__2483 (
            .O(N__10701),
            .I(N__10574));
    SRMux I__2482 (
            .O(N__10700),
            .I(N__10574));
    SRMux I__2481 (
            .O(N__10699),
            .I(N__10574));
    SRMux I__2480 (
            .O(N__10698),
            .I(N__10574));
    SRMux I__2479 (
            .O(N__10697),
            .I(N__10574));
    SRMux I__2478 (
            .O(N__10696),
            .I(N__10574));
    SRMux I__2477 (
            .O(N__10695),
            .I(N__10574));
    SRMux I__2476 (
            .O(N__10694),
            .I(N__10574));
    Glb2LocalMux I__2475 (
            .O(N__10691),
            .I(N__10574));
    SRMux I__2474 (
            .O(N__10690),
            .I(N__10574));
    SRMux I__2473 (
            .O(N__10689),
            .I(N__10574));
    SRMux I__2472 (
            .O(N__10688),
            .I(N__10574));
    SRMux I__2471 (
            .O(N__10687),
            .I(N__10574));
    SRMux I__2470 (
            .O(N__10686),
            .I(N__10574));
    Glb2LocalMux I__2469 (
            .O(N__10683),
            .I(N__10574));
    SRMux I__2468 (
            .O(N__10682),
            .I(N__10574));
    SRMux I__2467 (
            .O(N__10681),
            .I(N__10574));
    SRMux I__2466 (
            .O(N__10680),
            .I(N__10574));
    SRMux I__2465 (
            .O(N__10679),
            .I(N__10574));
    Glb2LocalMux I__2464 (
            .O(N__10676),
            .I(N__10574));
    SRMux I__2463 (
            .O(N__10675),
            .I(N__10574));
    SRMux I__2462 (
            .O(N__10674),
            .I(N__10574));
    SRMux I__2461 (
            .O(N__10673),
            .I(N__10574));
    SRMux I__2460 (
            .O(N__10672),
            .I(N__10574));
    SRMux I__2459 (
            .O(N__10671),
            .I(N__10574));
    SRMux I__2458 (
            .O(N__10670),
            .I(N__10574));
    SRMux I__2457 (
            .O(N__10669),
            .I(N__10574));
    SRMux I__2456 (
            .O(N__10668),
            .I(N__10574));
    SRMux I__2455 (
            .O(N__10667),
            .I(N__10574));
    SRMux I__2454 (
            .O(N__10666),
            .I(N__10574));
    SRMux I__2453 (
            .O(N__10665),
            .I(N__10574));
    SRMux I__2452 (
            .O(N__10664),
            .I(N__10574));
    SRMux I__2451 (
            .O(N__10663),
            .I(N__10574));
    SRMux I__2450 (
            .O(N__10662),
            .I(N__10574));
    SRMux I__2449 (
            .O(N__10661),
            .I(N__10574));
    Glb2LocalMux I__2448 (
            .O(N__10658),
            .I(N__10574));
    SRMux I__2447 (
            .O(N__10657),
            .I(N__10574));
    GlobalMux I__2446 (
            .O(N__10574),
            .I(N__10571));
    gio2CtrlBuf I__2445 (
            .O(N__10571),
            .I(RESETn_c_i_g));
    CascadeMux I__2444 (
            .O(N__10568),
            .I(N__10564));
    InMux I__2443 (
            .O(N__10567),
            .I(N__10555));
    InMux I__2442 (
            .O(N__10564),
            .I(N__10542));
    InMux I__2441 (
            .O(N__10563),
            .I(N__10535));
    InMux I__2440 (
            .O(N__10562),
            .I(N__10535));
    InMux I__2439 (
            .O(N__10561),
            .I(N__10535));
    InMux I__2438 (
            .O(N__10560),
            .I(N__10528));
    InMux I__2437 (
            .O(N__10559),
            .I(N__10528));
    InMux I__2436 (
            .O(N__10558),
            .I(N__10528));
    LocalMux I__2435 (
            .O(N__10555),
            .I(N__10525));
    InMux I__2434 (
            .O(N__10554),
            .I(N__10516));
    InMux I__2433 (
            .O(N__10553),
            .I(N__10516));
    InMux I__2432 (
            .O(N__10552),
            .I(N__10516));
    InMux I__2431 (
            .O(N__10551),
            .I(N__10516));
    InMux I__2430 (
            .O(N__10550),
            .I(N__10511));
    InMux I__2429 (
            .O(N__10549),
            .I(N__10511));
    InMux I__2428 (
            .O(N__10548),
            .I(N__10501));
    InMux I__2427 (
            .O(N__10547),
            .I(N__10496));
    InMux I__2426 (
            .O(N__10546),
            .I(N__10496));
    InMux I__2425 (
            .O(N__10545),
            .I(N__10493));
    LocalMux I__2424 (
            .O(N__10542),
            .I(N__10481));
    LocalMux I__2423 (
            .O(N__10535),
            .I(N__10481));
    LocalMux I__2422 (
            .O(N__10528),
            .I(N__10478));
    Span4Mux_v I__2421 (
            .O(N__10525),
            .I(N__10471));
    LocalMux I__2420 (
            .O(N__10516),
            .I(N__10471));
    LocalMux I__2419 (
            .O(N__10511),
            .I(N__10471));
    InMux I__2418 (
            .O(N__10510),
            .I(N__10464));
    InMux I__2417 (
            .O(N__10509),
            .I(N__10464));
    InMux I__2416 (
            .O(N__10508),
            .I(N__10453));
    InMux I__2415 (
            .O(N__10507),
            .I(N__10453));
    InMux I__2414 (
            .O(N__10506),
            .I(N__10453));
    InMux I__2413 (
            .O(N__10505),
            .I(N__10453));
    InMux I__2412 (
            .O(N__10504),
            .I(N__10453));
    LocalMux I__2411 (
            .O(N__10501),
            .I(N__10446));
    LocalMux I__2410 (
            .O(N__10496),
            .I(N__10446));
    LocalMux I__2409 (
            .O(N__10493),
            .I(N__10446));
    InMux I__2408 (
            .O(N__10492),
            .I(N__10439));
    InMux I__2407 (
            .O(N__10491),
            .I(N__10439));
    InMux I__2406 (
            .O(N__10490),
            .I(N__10439));
    InMux I__2405 (
            .O(N__10489),
            .I(N__10432));
    InMux I__2404 (
            .O(N__10488),
            .I(N__10432));
    InMux I__2403 (
            .O(N__10487),
            .I(N__10432));
    InMux I__2402 (
            .O(N__10486),
            .I(N__10429));
    Span4Mux_v I__2401 (
            .O(N__10481),
            .I(N__10417));
    Span4Mux_v I__2400 (
            .O(N__10478),
            .I(N__10417));
    Span4Mux_v I__2399 (
            .O(N__10471),
            .I(N__10417));
    InMux I__2398 (
            .O(N__10470),
            .I(N__10414));
    InMux I__2397 (
            .O(N__10469),
            .I(N__10409));
    LocalMux I__2396 (
            .O(N__10464),
            .I(N__10406));
    LocalMux I__2395 (
            .O(N__10453),
            .I(N__10395));
    Span4Mux_v I__2394 (
            .O(N__10446),
            .I(N__10395));
    LocalMux I__2393 (
            .O(N__10439),
            .I(N__10395));
    LocalMux I__2392 (
            .O(N__10432),
            .I(N__10395));
    LocalMux I__2391 (
            .O(N__10429),
            .I(N__10395));
    InMux I__2390 (
            .O(N__10428),
            .I(N__10390));
    InMux I__2389 (
            .O(N__10427),
            .I(N__10390));
    InMux I__2388 (
            .O(N__10426),
            .I(N__10383));
    InMux I__2387 (
            .O(N__10425),
            .I(N__10383));
    InMux I__2386 (
            .O(N__10424),
            .I(N__10383));
    Span4Mux_h I__2385 (
            .O(N__10417),
            .I(N__10380));
    LocalMux I__2384 (
            .O(N__10414),
            .I(N__10377));
    InMux I__2383 (
            .O(N__10413),
            .I(N__10372));
    InMux I__2382 (
            .O(N__10412),
            .I(N__10372));
    LocalMux I__2381 (
            .O(N__10409),
            .I(N__10369));
    Span4Mux_v I__2380 (
            .O(N__10406),
            .I(N__10364));
    Span4Mux_v I__2379 (
            .O(N__10395),
            .I(N__10364));
    LocalMux I__2378 (
            .O(N__10390),
            .I(N__10359));
    LocalMux I__2377 (
            .O(N__10383),
            .I(N__10359));
    Span4Mux_h I__2376 (
            .O(N__10380),
            .I(N__10354));
    Span4Mux_v I__2375 (
            .O(N__10377),
            .I(N__10354));
    LocalMux I__2374 (
            .O(N__10372),
            .I(N__10351));
    Span12Mux_v I__2373 (
            .O(N__10369),
            .I(N__10344));
    Sp12to4 I__2372 (
            .O(N__10364),
            .I(N__10344));
    Span12Mux_v I__2371 (
            .O(N__10359),
            .I(N__10344));
    Span4Mux_h I__2370 (
            .O(N__10354),
            .I(N__10341));
    Span12Mux_h I__2369 (
            .O(N__10351),
            .I(N__10338));
    Span12Mux_h I__2368 (
            .O(N__10344),
            .I(N__10335));
    Span4Mux_h I__2367 (
            .O(N__10341),
            .I(N__10332));
    Odrv12 I__2366 (
            .O(N__10338),
            .I(RESETn_c));
    Odrv12 I__2365 (
            .O(N__10335),
            .I(RESETn_c));
    Odrv4 I__2364 (
            .O(N__10332),
            .I(RESETn_c));
    InMux I__2363 (
            .O(N__10325),
            .I(N__10322));
    LocalMux I__2362 (
            .O(N__10322),
            .I(N__10319));
    Span12Mux_h I__2361 (
            .O(N__10319),
            .I(N__10316));
    Odrv12 I__2360 (
            .O(N__10316),
            .I(RAS1n_c));
    InMux I__2359 (
            .O(N__10313),
            .I(N__10310));
    LocalMux I__2358 (
            .O(N__10310),
            .I(N__10306));
    InMux I__2357 (
            .O(N__10309),
            .I(N__10303));
    Sp12to4 I__2356 (
            .O(N__10306),
            .I(N__10300));
    LocalMux I__2355 (
            .O(N__10303),
            .I(N__10297));
    Span12Mux_v I__2354 (
            .O(N__10300),
            .I(N__10294));
    Span12Mux_h I__2353 (
            .O(N__10297),
            .I(N__10291));
    Odrv12 I__2352 (
            .O(N__10294),
            .I(RAS0n_c));
    Odrv12 I__2351 (
            .O(N__10291),
            .I(RAS0n_c));
    InMux I__2350 (
            .O(N__10286),
            .I(N__10283));
    LocalMux I__2349 (
            .O(N__10283),
            .I(N__10280));
    Span12Mux_v I__2348 (
            .O(N__10280),
            .I(N__10277));
    Odrv12 I__2347 (
            .O(N__10277),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ));
    InMux I__2346 (
            .O(N__10274),
            .I(N__10271));
    LocalMux I__2345 (
            .O(N__10271),
            .I(N__10243));
    ClkMux I__2344 (
            .O(N__10270),
            .I(N__10136));
    ClkMux I__2343 (
            .O(N__10269),
            .I(N__10136));
    ClkMux I__2342 (
            .O(N__10268),
            .I(N__10136));
    ClkMux I__2341 (
            .O(N__10267),
            .I(N__10136));
    ClkMux I__2340 (
            .O(N__10266),
            .I(N__10136));
    ClkMux I__2339 (
            .O(N__10265),
            .I(N__10136));
    ClkMux I__2338 (
            .O(N__10264),
            .I(N__10136));
    ClkMux I__2337 (
            .O(N__10263),
            .I(N__10136));
    ClkMux I__2336 (
            .O(N__10262),
            .I(N__10136));
    ClkMux I__2335 (
            .O(N__10261),
            .I(N__10136));
    ClkMux I__2334 (
            .O(N__10260),
            .I(N__10136));
    ClkMux I__2333 (
            .O(N__10259),
            .I(N__10136));
    ClkMux I__2332 (
            .O(N__10258),
            .I(N__10136));
    ClkMux I__2331 (
            .O(N__10257),
            .I(N__10136));
    ClkMux I__2330 (
            .O(N__10256),
            .I(N__10136));
    ClkMux I__2329 (
            .O(N__10255),
            .I(N__10136));
    ClkMux I__2328 (
            .O(N__10254),
            .I(N__10136));
    ClkMux I__2327 (
            .O(N__10253),
            .I(N__10136));
    ClkMux I__2326 (
            .O(N__10252),
            .I(N__10136));
    ClkMux I__2325 (
            .O(N__10251),
            .I(N__10136));
    ClkMux I__2324 (
            .O(N__10250),
            .I(N__10136));
    ClkMux I__2323 (
            .O(N__10249),
            .I(N__10136));
    ClkMux I__2322 (
            .O(N__10248),
            .I(N__10136));
    ClkMux I__2321 (
            .O(N__10247),
            .I(N__10136));
    ClkMux I__2320 (
            .O(N__10246),
            .I(N__10136));
    Glb2LocalMux I__2319 (
            .O(N__10243),
            .I(N__10136));
    ClkMux I__2318 (
            .O(N__10242),
            .I(N__10136));
    ClkMux I__2317 (
            .O(N__10241),
            .I(N__10136));
    ClkMux I__2316 (
            .O(N__10240),
            .I(N__10136));
    ClkMux I__2315 (
            .O(N__10239),
            .I(N__10136));
    ClkMux I__2314 (
            .O(N__10238),
            .I(N__10136));
    ClkMux I__2313 (
            .O(N__10237),
            .I(N__10136));
    ClkMux I__2312 (
            .O(N__10236),
            .I(N__10136));
    ClkMux I__2311 (
            .O(N__10235),
            .I(N__10136));
    ClkMux I__2310 (
            .O(N__10234),
            .I(N__10136));
    ClkMux I__2309 (
            .O(N__10233),
            .I(N__10136));
    ClkMux I__2308 (
            .O(N__10232),
            .I(N__10136));
    ClkMux I__2307 (
            .O(N__10231),
            .I(N__10136));
    ClkMux I__2306 (
            .O(N__10230),
            .I(N__10136));
    ClkMux I__2305 (
            .O(N__10229),
            .I(N__10136));
    ClkMux I__2304 (
            .O(N__10228),
            .I(N__10136));
    ClkMux I__2303 (
            .O(N__10227),
            .I(N__10136));
    ClkMux I__2302 (
            .O(N__10226),
            .I(N__10136));
    ClkMux I__2301 (
            .O(N__10225),
            .I(N__10136));
    GlobalMux I__2300 (
            .O(N__10136),
            .I(CLK80_PLL));
    InMux I__2299 (
            .O(N__10133),
            .I(N__10130));
    LocalMux I__2298 (
            .O(N__10130),
            .I(N__10127));
    Span4Mux_v I__2297 (
            .O(N__10127),
            .I(N__10123));
    InMux I__2296 (
            .O(N__10126),
            .I(N__10120));
    Sp12to4 I__2295 (
            .O(N__10123),
            .I(N__10117));
    LocalMux I__2294 (
            .O(N__10120),
            .I(N__10114));
    Span12Mux_h I__2293 (
            .O(N__10117),
            .I(N__10107));
    Span12Mux_h I__2292 (
            .O(N__10114),
            .I(N__10107));
    InMux I__2291 (
            .O(N__10113),
            .I(N__10104));
    InMux I__2290 (
            .O(N__10112),
            .I(N__10101));
    Odrv12 I__2289 (
            .O(N__10107),
            .I(REG_CYCLEm));
    LocalMux I__2288 (
            .O(N__10104),
            .I(REG_CYCLEm));
    LocalMux I__2287 (
            .O(N__10101),
            .I(REG_CYCLEm));
    CascadeMux I__2286 (
            .O(N__10094),
            .I(N__10091));
    InMux I__2285 (
            .O(N__10091),
            .I(N__10086));
    CascadeMux I__2284 (
            .O(N__10090),
            .I(N__10083));
    CascadeMux I__2283 (
            .O(N__10089),
            .I(N__10080));
    LocalMux I__2282 (
            .O(N__10086),
            .I(N__10076));
    InMux I__2281 (
            .O(N__10083),
            .I(N__10071));
    InMux I__2280 (
            .O(N__10080),
            .I(N__10071));
    CascadeMux I__2279 (
            .O(N__10079),
            .I(N__10066));
    Span4Mux_v I__2278 (
            .O(N__10076),
            .I(N__10063));
    LocalMux I__2277 (
            .O(N__10071),
            .I(N__10060));
    InMux I__2276 (
            .O(N__10070),
            .I(N__10056));
    InMux I__2275 (
            .O(N__10069),
            .I(N__10053));
    InMux I__2274 (
            .O(N__10066),
            .I(N__10046));
    Sp12to4 I__2273 (
            .O(N__10063),
            .I(N__10043));
    Span4Mux_v I__2272 (
            .O(N__10060),
            .I(N__10038));
    InMux I__2271 (
            .O(N__10059),
            .I(N__10035));
    LocalMux I__2270 (
            .O(N__10056),
            .I(N__10030));
    LocalMux I__2269 (
            .O(N__10053),
            .I(N__10030));
    InMux I__2268 (
            .O(N__10052),
            .I(N__10025));
    InMux I__2267 (
            .O(N__10051),
            .I(N__10020));
    InMux I__2266 (
            .O(N__10050),
            .I(N__10020));
    InMux I__2265 (
            .O(N__10049),
            .I(N__10017));
    LocalMux I__2264 (
            .O(N__10046),
            .I(N__10013));
    Span12Mux_s9_h I__2263 (
            .O(N__10043),
            .I(N__10007));
    InMux I__2262 (
            .O(N__10042),
            .I(N__10002));
    InMux I__2261 (
            .O(N__10041),
            .I(N__10002));
    Span4Mux_h I__2260 (
            .O(N__10038),
            .I(N__9994));
    LocalMux I__2259 (
            .O(N__10035),
            .I(N__9994));
    Span4Mux_v I__2258 (
            .O(N__10030),
            .I(N__9989));
    InMux I__2257 (
            .O(N__10029),
            .I(N__9984));
    InMux I__2256 (
            .O(N__10028),
            .I(N__9984));
    LocalMux I__2255 (
            .O(N__10025),
            .I(N__9977));
    LocalMux I__2254 (
            .O(N__10020),
            .I(N__9977));
    LocalMux I__2253 (
            .O(N__10017),
            .I(N__9977));
    InMux I__2252 (
            .O(N__10016),
            .I(N__9974));
    Span4Mux_h I__2251 (
            .O(N__10013),
            .I(N__9971));
    InMux I__2250 (
            .O(N__10012),
            .I(N__9964));
    InMux I__2249 (
            .O(N__10011),
            .I(N__9964));
    InMux I__2248 (
            .O(N__10010),
            .I(N__9964));
    Span12Mux_v I__2247 (
            .O(N__10007),
            .I(N__9959));
    LocalMux I__2246 (
            .O(N__10002),
            .I(N__9959));
    InMux I__2245 (
            .O(N__10001),
            .I(N__9952));
    InMux I__2244 (
            .O(N__10000),
            .I(N__9952));
    InMux I__2243 (
            .O(N__9999),
            .I(N__9952));
    Span4Mux_v I__2242 (
            .O(N__9994),
            .I(N__9949));
    InMux I__2241 (
            .O(N__9993),
            .I(N__9944));
    InMux I__2240 (
            .O(N__9992),
            .I(N__9944));
    Span4Mux_v I__2239 (
            .O(N__9989),
            .I(N__9937));
    LocalMux I__2238 (
            .O(N__9984),
            .I(N__9937));
    Span4Mux_v I__2237 (
            .O(N__9977),
            .I(N__9937));
    LocalMux I__2236 (
            .O(N__9974),
            .I(N__9934));
    Odrv4 I__2235 (
            .O(N__9971),
            .I(CPU_CYCLEm));
    LocalMux I__2234 (
            .O(N__9964),
            .I(CPU_CYCLEm));
    Odrv12 I__2233 (
            .O(N__9959),
            .I(CPU_CYCLEm));
    LocalMux I__2232 (
            .O(N__9952),
            .I(CPU_CYCLEm));
    Odrv4 I__2231 (
            .O(N__9949),
            .I(CPU_CYCLEm));
    LocalMux I__2230 (
            .O(N__9944),
            .I(CPU_CYCLEm));
    Odrv4 I__2229 (
            .O(N__9937),
            .I(CPU_CYCLEm));
    Odrv4 I__2228 (
            .O(N__9934),
            .I(CPU_CYCLEm));
    IoInMux I__2227 (
            .O(N__9917),
            .I(N__9914));
    LocalMux I__2226 (
            .O(N__9914),
            .I(N__9911));
    Span4Mux_s3_v I__2225 (
            .O(N__9911),
            .I(N__9908));
    Span4Mux_v I__2224 (
            .O(N__9908),
            .I(N__9905));
    Odrv4 I__2223 (
            .O(N__9905),
            .I(N_136_i));
    CascadeMux I__2222 (
            .O(N__9902),
            .I(N__9898));
    InMux I__2221 (
            .O(N__9901),
            .I(N__9895));
    InMux I__2220 (
            .O(N__9898),
            .I(N__9891));
    LocalMux I__2219 (
            .O(N__9895),
            .I(N__9888));
    InMux I__2218 (
            .O(N__9894),
            .I(N__9885));
    LocalMux I__2217 (
            .O(N__9891),
            .I(N__9882));
    Span4Mux_v I__2216 (
            .O(N__9888),
            .I(N__9879));
    LocalMux I__2215 (
            .O(N__9885),
            .I(N__9876));
    Span4Mux_v I__2214 (
            .O(N__9882),
            .I(N__9872));
    Span4Mux_v I__2213 (
            .O(N__9879),
            .I(N__9867));
    Span4Mux_h I__2212 (
            .O(N__9876),
            .I(N__9867));
    CascadeMux I__2211 (
            .O(N__9875),
            .I(N__9864));
    Span4Mux_v I__2210 (
            .O(N__9872),
            .I(N__9859));
    Span4Mux_h I__2209 (
            .O(N__9867),
            .I(N__9859));
    InMux I__2208 (
            .O(N__9864),
            .I(N__9854));
    Span4Mux_h I__2207 (
            .O(N__9859),
            .I(N__9851));
    InMux I__2206 (
            .O(N__9858),
            .I(N__9846));
    InMux I__2205 (
            .O(N__9857),
            .I(N__9846));
    LocalMux I__2204 (
            .O(N__9854),
            .I(N__9843));
    Span4Mux_h I__2203 (
            .O(N__9851),
            .I(N__9838));
    LocalMux I__2202 (
            .O(N__9846),
            .I(N__9838));
    Span12Mux_v I__2201 (
            .O(N__9843),
            .I(N__9835));
    Span4Mux_h I__2200 (
            .O(N__9838),
            .I(N__9832));
    Span12Mux_h I__2199 (
            .O(N__9835),
            .I(N__9829));
    Span4Mux_v I__2198 (
            .O(N__9832),
            .I(N__9826));
    Odrv12 I__2197 (
            .O(N__9829),
            .I(CASUn_c));
    Odrv4 I__2196 (
            .O(N__9826),
            .I(CASUn_c));
    InMux I__2195 (
            .O(N__9821),
            .I(N__9817));
    InMux I__2194 (
            .O(N__9820),
            .I(N__9814));
    LocalMux I__2193 (
            .O(N__9817),
            .I(N__9811));
    LocalMux I__2192 (
            .O(N__9814),
            .I(N__9805));
    Span4Mux_v I__2191 (
            .O(N__9811),
            .I(N__9802));
    InMux I__2190 (
            .O(N__9810),
            .I(N__9799));
    CascadeMux I__2189 (
            .O(N__9809),
            .I(N__9796));
    InMux I__2188 (
            .O(N__9808),
            .I(N__9793));
    Span4Mux_v I__2187 (
            .O(N__9805),
            .I(N__9790));
    Span4Mux_v I__2186 (
            .O(N__9802),
            .I(N__9785));
    LocalMux I__2185 (
            .O(N__9799),
            .I(N__9785));
    InMux I__2184 (
            .O(N__9796),
            .I(N__9782));
    LocalMux I__2183 (
            .O(N__9793),
            .I(N__9779));
    Sp12to4 I__2182 (
            .O(N__9790),
            .I(N__9776));
    Span4Mux_v I__2181 (
            .O(N__9785),
            .I(N__9773));
    LocalMux I__2180 (
            .O(N__9782),
            .I(N__9768));
    Sp12to4 I__2179 (
            .O(N__9779),
            .I(N__9768));
    Span12Mux_h I__2178 (
            .O(N__9776),
            .I(N__9763));
    Sp12to4 I__2177 (
            .O(N__9773),
            .I(N__9763));
    Span12Mux_v I__2176 (
            .O(N__9768),
            .I(N__9760));
    Span12Mux_h I__2175 (
            .O(N__9763),
            .I(N__9757));
    Span12Mux_h I__2174 (
            .O(N__9760),
            .I(N__9754));
    Odrv12 I__2173 (
            .O(N__9757),
            .I(RnW_c));
    Odrv12 I__2172 (
            .O(N__9754),
            .I(RnW_c));
    InMux I__2171 (
            .O(N__9749),
            .I(N__9741));
    InMux I__2170 (
            .O(N__9748),
            .I(N__9741));
    InMux I__2169 (
            .O(N__9747),
            .I(N__9736));
    InMux I__2168 (
            .O(N__9746),
            .I(N__9736));
    LocalMux I__2167 (
            .O(N__9741),
            .I(N__9733));
    LocalMux I__2166 (
            .O(N__9736),
            .I(N__9730));
    Span4Mux_v I__2165 (
            .O(N__9733),
            .I(N__9727));
    Span4Mux_v I__2164 (
            .O(N__9730),
            .I(N__9724));
    Sp12to4 I__2163 (
            .O(N__9727),
            .I(N__9721));
    Span4Mux_h I__2162 (
            .O(N__9724),
            .I(N__9718));
    Span12Mux_h I__2161 (
            .O(N__9721),
            .I(N__9713));
    Sp12to4 I__2160 (
            .O(N__9718),
            .I(N__9713));
    Odrv12 I__2159 (
            .O(N__9713),
            .I(DRA_c_7));
    InMux I__2158 (
            .O(N__9710),
            .I(N__9705));
    InMux I__2157 (
            .O(N__9709),
            .I(N__9700));
    InMux I__2156 (
            .O(N__9708),
            .I(N__9700));
    LocalMux I__2155 (
            .O(N__9705),
            .I(N__9694));
    LocalMux I__2154 (
            .O(N__9700),
            .I(N__9694));
    InMux I__2153 (
            .O(N__9699),
            .I(N__9691));
    Sp12to4 I__2152 (
            .O(N__9694),
            .I(N__9686));
    LocalMux I__2151 (
            .O(N__9691),
            .I(N__9686));
    Span12Mux_v I__2150 (
            .O(N__9686),
            .I(N__9683));
    Span12Mux_h I__2149 (
            .O(N__9683),
            .I(N__9680));
    Odrv12 I__2148 (
            .O(N__9680),
            .I(DRA_c_6));
    InMux I__2147 (
            .O(N__9677),
            .I(N__9674));
    LocalMux I__2146 (
            .O(N__9674),
            .I(N__9671));
    Odrv4 I__2145 (
            .O(N__9671),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ));
    InMux I__2144 (
            .O(N__9668),
            .I(N__9665));
    LocalMux I__2143 (
            .O(N__9665),
            .I(N__9662));
    Span4Mux_h I__2142 (
            .O(N__9662),
            .I(N__9659));
    Odrv4 I__2141 (
            .O(N__9659),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ));
    InMux I__2140 (
            .O(N__9656),
            .I(N__9652));
    InMux I__2139 (
            .O(N__9655),
            .I(N__9647));
    LocalMux I__2138 (
            .O(N__9652),
            .I(N__9644));
    InMux I__2137 (
            .O(N__9651),
            .I(N__9641));
    InMux I__2136 (
            .O(N__9650),
            .I(N__9638));
    LocalMux I__2135 (
            .O(N__9647),
            .I(N__9635));
    Span4Mux_h I__2134 (
            .O(N__9644),
            .I(N__9628));
    LocalMux I__2133 (
            .O(N__9641),
            .I(N__9628));
    LocalMux I__2132 (
            .O(N__9638),
            .I(N__9628));
    Span4Mux_v I__2131 (
            .O(N__9635),
            .I(N__9625));
    Span4Mux_v I__2130 (
            .O(N__9628),
            .I(N__9622));
    Sp12to4 I__2129 (
            .O(N__9625),
            .I(N__9619));
    Span4Mux_v I__2128 (
            .O(N__9622),
            .I(N__9616));
    Span12Mux_h I__2127 (
            .O(N__9619),
            .I(N__9613));
    Sp12to4 I__2126 (
            .O(N__9616),
            .I(N__9610));
    Span12Mux_v I__2125 (
            .O(N__9613),
            .I(N__9607));
    Span12Mux_h I__2124 (
            .O(N__9610),
            .I(N__9604));
    Odrv12 I__2123 (
            .O(N__9607),
            .I(DRA_c_4));
    Odrv12 I__2122 (
            .O(N__9604),
            .I(DRA_c_4));
    InMux I__2121 (
            .O(N__9599),
            .I(N__9596));
    LocalMux I__2120 (
            .O(N__9596),
            .I(N__9590));
    InMux I__2119 (
            .O(N__9595),
            .I(N__9587));
    InMux I__2118 (
            .O(N__9594),
            .I(N__9584));
    InMux I__2117 (
            .O(N__9593),
            .I(N__9581));
    Sp12to4 I__2116 (
            .O(N__9590),
            .I(N__9572));
    LocalMux I__2115 (
            .O(N__9587),
            .I(N__9572));
    LocalMux I__2114 (
            .O(N__9584),
            .I(N__9572));
    LocalMux I__2113 (
            .O(N__9581),
            .I(N__9572));
    Span12Mux_v I__2112 (
            .O(N__9572),
            .I(N__9569));
    Span12Mux_h I__2111 (
            .O(N__9569),
            .I(N__9566));
    Odrv12 I__2110 (
            .O(N__9566),
            .I(DRA_c_3));
    InMux I__2109 (
            .O(N__9563),
            .I(N__9560));
    LocalMux I__2108 (
            .O(N__9560),
            .I(N__9557));
    Span4Mux_h I__2107 (
            .O(N__9557),
            .I(N__9554));
    Odrv4 I__2106 (
            .O(N__9554),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ));
    IoInMux I__2105 (
            .O(N__9551),
            .I(N__9548));
    LocalMux I__2104 (
            .O(N__9548),
            .I(N__9545));
    Span4Mux_s2_h I__2103 (
            .O(N__9545),
            .I(N__9542));
    Sp12to4 I__2102 (
            .O(N__9542),
            .I(N__9539));
    Span12Mux_v I__2101 (
            .O(N__9539),
            .I(N__9536));
    Span12Mux_h I__2100 (
            .O(N__9536),
            .I(N__9533));
    Odrv12 I__2099 (
            .O(N__9533),
            .I(N_146_i));
    CascadeMux I__2098 (
            .O(N__9530),
            .I(N__9524));
    InMux I__2097 (
            .O(N__9529),
            .I(N__9521));
    InMux I__2096 (
            .O(N__9528),
            .I(N__9516));
    InMux I__2095 (
            .O(N__9527),
            .I(N__9516));
    InMux I__2094 (
            .O(N__9524),
            .I(N__9513));
    LocalMux I__2093 (
            .O(N__9521),
            .I(N__9510));
    LocalMux I__2092 (
            .O(N__9516),
            .I(N__9505));
    LocalMux I__2091 (
            .O(N__9513),
            .I(N__9505));
    Span4Mux_v I__2090 (
            .O(N__9510),
            .I(N__9502));
    Span4Mux_v I__2089 (
            .O(N__9505),
            .I(N__9499));
    Sp12to4 I__2088 (
            .O(N__9502),
            .I(N__9496));
    Span4Mux_h I__2087 (
            .O(N__9499),
            .I(N__9493));
    Span12Mux_h I__2086 (
            .O(N__9496),
            .I(N__9488));
    Sp12to4 I__2085 (
            .O(N__9493),
            .I(N__9488));
    Span12Mux_v I__2084 (
            .O(N__9488),
            .I(N__9485));
    Odrv12 I__2083 (
            .O(N__9485),
            .I(CLK40_PLL_i));
    IoInMux I__2082 (
            .O(N__9482),
            .I(N__9478));
    IoInMux I__2081 (
            .O(N__9481),
            .I(N__9475));
    LocalMux I__2080 (
            .O(N__9478),
            .I(N__9472));
    LocalMux I__2079 (
            .O(N__9475),
            .I(N__9468));
    Span4Mux_s2_v I__2078 (
            .O(N__9472),
            .I(N__9465));
    IoInMux I__2077 (
            .O(N__9471),
            .I(N__9462));
    IoSpan4Mux I__2076 (
            .O(N__9468),
            .I(N__9459));
    Sp12to4 I__2075 (
            .O(N__9465),
            .I(N__9456));
    LocalMux I__2074 (
            .O(N__9462),
            .I(N__9453));
    Span4Mux_s2_h I__2073 (
            .O(N__9459),
            .I(N__9450));
    Span12Mux_h I__2072 (
            .O(N__9456),
            .I(N__9447));
    Span12Mux_s2_v I__2071 (
            .O(N__9453),
            .I(N__9444));
    Sp12to4 I__2070 (
            .O(N__9450),
            .I(N__9441));
    Span12Mux_v I__2069 (
            .O(N__9447),
            .I(N__9436));
    Span12Mux_v I__2068 (
            .O(N__9444),
            .I(N__9436));
    Span12Mux_s8_h I__2067 (
            .O(N__9441),
            .I(N__9433));
    Odrv12 I__2066 (
            .O(N__9436),
            .I(CLK40_PLL_i_i));
    Odrv12 I__2065 (
            .O(N__9433),
            .I(CLK40_PLL_i_i));
    InMux I__2064 (
            .O(N__9428),
            .I(N__9425));
    LocalMux I__2063 (
            .O(N__9425),
            .I(\U712_BYTE_ENABLE.N_406 ));
    InMux I__2062 (
            .O(N__9422),
            .I(N__9416));
    InMux I__2061 (
            .O(N__9421),
            .I(N__9416));
    LocalMux I__2060 (
            .O(N__9416),
            .I(\U712_BYTE_ENABLE.N_284_i ));
    IoInMux I__2059 (
            .O(N__9413),
            .I(N__9410));
    LocalMux I__2058 (
            .O(N__9410),
            .I(N__9407));
    IoSpan4Mux I__2057 (
            .O(N__9407),
            .I(N__9404));
    Span4Mux_s2_v I__2056 (
            .O(N__9404),
            .I(N__9401));
    Span4Mux_v I__2055 (
            .O(N__9401),
            .I(N__9398));
    Odrv4 I__2054 (
            .O(N__9398),
            .I(N_374_i));
    CascadeMux I__2053 (
            .O(N__9395),
            .I(N__9392));
    InMux I__2052 (
            .O(N__9392),
            .I(N__9388));
    InMux I__2051 (
            .O(N__9391),
            .I(N__9385));
    LocalMux I__2050 (
            .O(N__9388),
            .I(\U712_BYTE_ENABLE.N_409 ));
    LocalMux I__2049 (
            .O(N__9385),
            .I(\U712_BYTE_ENABLE.N_409 ));
    CascadeMux I__2048 (
            .O(N__9380),
            .I(N__9374));
    CascadeMux I__2047 (
            .O(N__9379),
            .I(N__9371));
    CascadeMux I__2046 (
            .O(N__9378),
            .I(N__9366));
    InMux I__2045 (
            .O(N__9377),
            .I(N__9356));
    InMux I__2044 (
            .O(N__9374),
            .I(N__9356));
    InMux I__2043 (
            .O(N__9371),
            .I(N__9356));
    InMux I__2042 (
            .O(N__9370),
            .I(N__9353));
    InMux I__2041 (
            .O(N__9369),
            .I(N__9349));
    InMux I__2040 (
            .O(N__9366),
            .I(N__9346));
    CascadeMux I__2039 (
            .O(N__9365),
            .I(N__9342));
    InMux I__2038 (
            .O(N__9364),
            .I(N__9339));
    InMux I__2037 (
            .O(N__9363),
            .I(N__9336));
    LocalMux I__2036 (
            .O(N__9356),
            .I(N__9331));
    LocalMux I__2035 (
            .O(N__9353),
            .I(N__9331));
    CascadeMux I__2034 (
            .O(N__9352),
            .I(N__9328));
    LocalMux I__2033 (
            .O(N__9349),
            .I(N__9322));
    LocalMux I__2032 (
            .O(N__9346),
            .I(N__9319));
    InMux I__2031 (
            .O(N__9345),
            .I(N__9316));
    InMux I__2030 (
            .O(N__9342),
            .I(N__9313));
    LocalMux I__2029 (
            .O(N__9339),
            .I(N__9310));
    LocalMux I__2028 (
            .O(N__9336),
            .I(N__9307));
    Span4Mux_h I__2027 (
            .O(N__9331),
            .I(N__9304));
    InMux I__2026 (
            .O(N__9328),
            .I(N__9301));
    InMux I__2025 (
            .O(N__9327),
            .I(N__9298));
    InMux I__2024 (
            .O(N__9326),
            .I(N__9295));
    InMux I__2023 (
            .O(N__9325),
            .I(N__9292));
    Span4Mux_v I__2022 (
            .O(N__9322),
            .I(N__9285));
    Span4Mux_v I__2021 (
            .O(N__9319),
            .I(N__9285));
    LocalMux I__2020 (
            .O(N__9316),
            .I(N__9285));
    LocalMux I__2019 (
            .O(N__9313),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2018 (
            .O(N__9310),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv12 I__2017 (
            .O(N__9307),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2016 (
            .O(N__9304),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2015 (
            .O(N__9301),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2014 (
            .O(N__9298),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2013 (
            .O(N__9295),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    LocalMux I__2012 (
            .O(N__9292),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    Odrv4 I__2011 (
            .O(N__9285),
            .I(\U712_REG_SM.C1_SYNCZ0Z_1 ));
    IoInMux I__2010 (
            .O(N__9266),
            .I(N__9263));
    LocalMux I__2009 (
            .O(N__9263),
            .I(N__9260));
    Span12Mux_s4_v I__2008 (
            .O(N__9260),
            .I(N__9257));
    Span12Mux_h I__2007 (
            .O(N__9257),
            .I(N__9254));
    Odrv12 I__2006 (
            .O(N__9254),
            .I(ASn_c));
    CEMux I__2005 (
            .O(N__9251),
            .I(N__9248));
    LocalMux I__2004 (
            .O(N__9248),
            .I(N__9245));
    Odrv4 I__2003 (
            .O(N__9245),
            .I(\U712_REG_SM.N_95_0 ));
    IoInMux I__2002 (
            .O(N__9242),
            .I(N__9239));
    LocalMux I__2001 (
            .O(N__9239),
            .I(N__9236));
    Span4Mux_s2_v I__2000 (
            .O(N__9236),
            .I(N__9233));
    Span4Mux_v I__1999 (
            .O(N__9233),
            .I(N__9230));
    Odrv4 I__1998 (
            .O(N__9230),
            .I(LLBEn_c));
    InMux I__1997 (
            .O(N__9227),
            .I(N__9221));
    CascadeMux I__1996 (
            .O(N__9226),
            .I(N__9211));
    CascadeMux I__1995 (
            .O(N__9225),
            .I(N__9206));
    InMux I__1994 (
            .O(N__9224),
            .I(N__9203));
    LocalMux I__1993 (
            .O(N__9221),
            .I(N__9200));
    InMux I__1992 (
            .O(N__9220),
            .I(N__9197));
    InMux I__1991 (
            .O(N__9219),
            .I(N__9186));
    InMux I__1990 (
            .O(N__9218),
            .I(N__9186));
    InMux I__1989 (
            .O(N__9217),
            .I(N__9186));
    InMux I__1988 (
            .O(N__9216),
            .I(N__9186));
    InMux I__1987 (
            .O(N__9215),
            .I(N__9186));
    InMux I__1986 (
            .O(N__9214),
            .I(N__9183));
    InMux I__1985 (
            .O(N__9211),
            .I(N__9180));
    CascadeMux I__1984 (
            .O(N__9210),
            .I(N__9177));
    CascadeMux I__1983 (
            .O(N__9209),
            .I(N__9174));
    InMux I__1982 (
            .O(N__9206),
            .I(N__9170));
    LocalMux I__1981 (
            .O(N__9203),
            .I(N__9153));
    Span4Mux_h I__1980 (
            .O(N__9200),
            .I(N__9153));
    LocalMux I__1979 (
            .O(N__9197),
            .I(N__9153));
    LocalMux I__1978 (
            .O(N__9186),
            .I(N__9153));
    LocalMux I__1977 (
            .O(N__9183),
            .I(N__9145));
    LocalMux I__1976 (
            .O(N__9180),
            .I(N__9145));
    InMux I__1975 (
            .O(N__9177),
            .I(N__9138));
    InMux I__1974 (
            .O(N__9174),
            .I(N__9138));
    InMux I__1973 (
            .O(N__9173),
            .I(N__9138));
    LocalMux I__1972 (
            .O(N__9170),
            .I(N__9134));
    InMux I__1971 (
            .O(N__9169),
            .I(N__9125));
    InMux I__1970 (
            .O(N__9168),
            .I(N__9125));
    InMux I__1969 (
            .O(N__9167),
            .I(N__9125));
    InMux I__1968 (
            .O(N__9166),
            .I(N__9125));
    InMux I__1967 (
            .O(N__9165),
            .I(N__9116));
    InMux I__1966 (
            .O(N__9164),
            .I(N__9116));
    InMux I__1965 (
            .O(N__9163),
            .I(N__9116));
    InMux I__1964 (
            .O(N__9162),
            .I(N__9116));
    Span4Mux_h I__1963 (
            .O(N__9153),
            .I(N__9113));
    InMux I__1962 (
            .O(N__9152),
            .I(N__9106));
    InMux I__1961 (
            .O(N__9151),
            .I(N__9106));
    InMux I__1960 (
            .O(N__9150),
            .I(N__9106));
    Span4Mux_h I__1959 (
            .O(N__9145),
            .I(N__9101));
    LocalMux I__1958 (
            .O(N__9138),
            .I(N__9101));
    InMux I__1957 (
            .O(N__9137),
            .I(N__9098));
    Odrv4 I__1956 (
            .O(N__9134),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1955 (
            .O(N__9125),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1954 (
            .O(N__9116),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1953 (
            .O(N__9113),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1952 (
            .O(N__9106),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    Odrv4 I__1951 (
            .O(N__9101),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    LocalMux I__1950 (
            .O(N__9098),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ));
    IoInMux I__1949 (
            .O(N__9083),
            .I(N__9080));
    LocalMux I__1948 (
            .O(N__9080),
            .I(N__9077));
    Span4Mux_s3_v I__1947 (
            .O(N__9077),
            .I(N__9074));
    Sp12to4 I__1946 (
            .O(N__9074),
            .I(N__9071));
    Span12Mux_h I__1945 (
            .O(N__9071),
            .I(N__9068));
    Odrv12 I__1944 (
            .O(N__9068),
            .I(CASn_c));
    InMux I__1943 (
            .O(N__9065),
            .I(N__9059));
    InMux I__1942 (
            .O(N__9064),
            .I(N__9056));
    InMux I__1941 (
            .O(N__9063),
            .I(N__9051));
    InMux I__1940 (
            .O(N__9062),
            .I(N__9051));
    LocalMux I__1939 (
            .O(N__9059),
            .I(N__9044));
    LocalMux I__1938 (
            .O(N__9056),
            .I(N__9044));
    LocalMux I__1937 (
            .O(N__9051),
            .I(N__9044));
    Sp12to4 I__1936 (
            .O(N__9044),
            .I(N__9041));
    Span12Mux_v I__1935 (
            .O(N__9041),
            .I(N__9038));
    Span12Mux_h I__1934 (
            .O(N__9038),
            .I(N__9035));
    Odrv12 I__1933 (
            .O(N__9035),
            .I(DRA_c_5));
    InMux I__1932 (
            .O(N__9032),
            .I(N__9029));
    LocalMux I__1931 (
            .O(N__9029),
            .I(N__9026));
    Odrv12 I__1930 (
            .O(N__9026),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ));
    InMux I__1929 (
            .O(N__9023),
            .I(N__9017));
    InMux I__1928 (
            .O(N__9022),
            .I(N__9017));
    LocalMux I__1927 (
            .O(N__9017),
            .I(N__9013));
    InMux I__1926 (
            .O(N__9016),
            .I(N__9010));
    Span4Mux_h I__1925 (
            .O(N__9013),
            .I(N__9004));
    LocalMux I__1924 (
            .O(N__9010),
            .I(N__9004));
    InMux I__1923 (
            .O(N__9009),
            .I(N__9001));
    Span4Mux_h I__1922 (
            .O(N__9004),
            .I(N__8996));
    LocalMux I__1921 (
            .O(N__9001),
            .I(N__8996));
    Sp12to4 I__1920 (
            .O(N__8996),
            .I(N__8993));
    Span12Mux_v I__1919 (
            .O(N__8993),
            .I(N__8990));
    Span12Mux_h I__1918 (
            .O(N__8990),
            .I(N__8987));
    Odrv12 I__1917 (
            .O(N__8987),
            .I(DRA_c_2));
    CascadeMux I__1916 (
            .O(N__8984),
            .I(N__8981));
    InMux I__1915 (
            .O(N__8981),
            .I(N__8978));
    LocalMux I__1914 (
            .O(N__8978),
            .I(N__8975));
    Span4Mux_v I__1913 (
            .O(N__8975),
            .I(N__8972));
    Odrv4 I__1912 (
            .O(N__8972),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ));
    CascadeMux I__1911 (
            .O(N__8969),
            .I(N__8964));
    InMux I__1910 (
            .O(N__8968),
            .I(N__8959));
    InMux I__1909 (
            .O(N__8967),
            .I(N__8959));
    InMux I__1908 (
            .O(N__8964),
            .I(N__8956));
    LocalMux I__1907 (
            .O(N__8959),
            .I(N__8952));
    LocalMux I__1906 (
            .O(N__8956),
            .I(N__8949));
    InMux I__1905 (
            .O(N__8955),
            .I(N__8946));
    Span4Mux_h I__1904 (
            .O(N__8952),
            .I(N__8939));
    Span4Mux_v I__1903 (
            .O(N__8949),
            .I(N__8939));
    LocalMux I__1902 (
            .O(N__8946),
            .I(N__8939));
    Span4Mux_h I__1901 (
            .O(N__8939),
            .I(N__8936));
    Sp12to4 I__1900 (
            .O(N__8936),
            .I(N__8933));
    Span12Mux_v I__1899 (
            .O(N__8933),
            .I(N__8930));
    Odrv12 I__1898 (
            .O(N__8930),
            .I(DRA_c_1));
    InMux I__1897 (
            .O(N__8927),
            .I(N__8923));
    InMux I__1896 (
            .O(N__8926),
            .I(N__8920));
    LocalMux I__1895 (
            .O(N__8923),
            .I(N__8917));
    LocalMux I__1894 (
            .O(N__8920),
            .I(N__8914));
    Span4Mux_v I__1893 (
            .O(N__8917),
            .I(N__8911));
    Span4Mux_v I__1892 (
            .O(N__8914),
            .I(N__8908));
    Sp12to4 I__1891 (
            .O(N__8911),
            .I(N__8905));
    Sp12to4 I__1890 (
            .O(N__8908),
            .I(N__8902));
    Span12Mux_h I__1889 (
            .O(N__8905),
            .I(N__8899));
    Span12Mux_h I__1888 (
            .O(N__8902),
            .I(N__8896));
    Span12Mux_v I__1887 (
            .O(N__8899),
            .I(N__8893));
    Span12Mux_v I__1886 (
            .O(N__8896),
            .I(N__8890));
    Odrv12 I__1885 (
            .O(N__8893),
            .I(DRA_c_0));
    Odrv12 I__1884 (
            .O(N__8890),
            .I(DRA_c_0));
    InMux I__1883 (
            .O(N__8885),
            .I(N__8882));
    LocalMux I__1882 (
            .O(N__8882),
            .I(N__8879));
    Span4Mux_v I__1881 (
            .O(N__8879),
            .I(N__8876));
    Odrv4 I__1880 (
            .O(N__8876),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ));
    InMux I__1879 (
            .O(N__8873),
            .I(N__8868));
    InMux I__1878 (
            .O(N__8872),
            .I(N__8865));
    InMux I__1877 (
            .O(N__8871),
            .I(N__8862));
    LocalMux I__1876 (
            .O(N__8868),
            .I(N__8857));
    LocalMux I__1875 (
            .O(N__8865),
            .I(N__8857));
    LocalMux I__1874 (
            .O(N__8862),
            .I(N__8854));
    Span4Mux_v I__1873 (
            .O(N__8857),
            .I(N__8850));
    Span4Mux_v I__1872 (
            .O(N__8854),
            .I(N__8847));
    InMux I__1871 (
            .O(N__8853),
            .I(N__8844));
    Sp12to4 I__1870 (
            .O(N__8850),
            .I(N__8837));
    Sp12to4 I__1869 (
            .O(N__8847),
            .I(N__8837));
    LocalMux I__1868 (
            .O(N__8844),
            .I(N__8837));
    Span12Mux_h I__1867 (
            .O(N__8837),
            .I(N__8834));
    Odrv12 I__1866 (
            .O(N__8834),
            .I(DRA_c_8));
    InMux I__1865 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__1864 (
            .O(N__8828),
            .I(N__8825));
    Odrv12 I__1863 (
            .O(N__8825),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ));
    InMux I__1862 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__1861 (
            .O(N__8819),
            .I(N__8816));
    Span4Mux_h I__1860 (
            .O(N__8816),
            .I(N__8813));
    Odrv4 I__1859 (
            .O(N__8813),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ));
    InMux I__1858 (
            .O(N__8810),
            .I(N__8807));
    LocalMux I__1857 (
            .O(N__8807),
            .I(N__8804));
    Odrv4 I__1856 (
            .O(N__8804),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ));
    InMux I__1855 (
            .O(N__8801),
            .I(N__8798));
    LocalMux I__1854 (
            .O(N__8798),
            .I(N__8795));
    Odrv4 I__1853 (
            .O(N__8795),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ));
    InMux I__1852 (
            .O(N__8792),
            .I(N__8789));
    LocalMux I__1851 (
            .O(N__8789),
            .I(N__8786));
    Span4Mux_h I__1850 (
            .O(N__8786),
            .I(N__8783));
    Odrv4 I__1849 (
            .O(N__8783),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ));
    InMux I__1848 (
            .O(N__8780),
            .I(N__8777));
    LocalMux I__1847 (
            .O(N__8777),
            .I(N__8774));
    Span4Mux_h I__1846 (
            .O(N__8774),
            .I(N__8771));
    Odrv4 I__1845 (
            .O(N__8771),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ));
    InMux I__1844 (
            .O(N__8768),
            .I(N__8762));
    InMux I__1843 (
            .O(N__8767),
            .I(N__8762));
    LocalMux I__1842 (
            .O(N__8762),
            .I(N__8759));
    Span4Mux_h I__1841 (
            .O(N__8759),
            .I(N__8756));
    Odrv4 I__1840 (
            .O(N__8756),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ));
    InMux I__1839 (
            .O(N__8753),
            .I(N__8750));
    LocalMux I__1838 (
            .O(N__8750),
            .I(N__8747));
    Span4Mux_v I__1837 (
            .O(N__8747),
            .I(N__8744));
    Odrv4 I__1836 (
            .O(N__8744),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ));
    InMux I__1835 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__1834 (
            .O(N__8738),
            .I(N__8735));
    Span4Mux_h I__1833 (
            .O(N__8735),
            .I(N__8732));
    Odrv4 I__1832 (
            .O(N__8732),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ));
    InMux I__1831 (
            .O(N__8729),
            .I(N__8726));
    LocalMux I__1830 (
            .O(N__8726),
            .I(N__8722));
    InMux I__1829 (
            .O(N__8725),
            .I(N__8719));
    Span4Mux_h I__1828 (
            .O(N__8722),
            .I(N__8716));
    LocalMux I__1827 (
            .O(N__8719),
            .I(N__8713));
    Span4Mux_v I__1826 (
            .O(N__8716),
            .I(N__8710));
    Span4Mux_v I__1825 (
            .O(N__8713),
            .I(N__8707));
    Odrv4 I__1824 (
            .O(N__8710),
            .I(DBRn_c_i));
    Odrv4 I__1823 (
            .O(N__8707),
            .I(DBRn_c_i));
    InMux I__1822 (
            .O(N__8702),
            .I(N__8699));
    LocalMux I__1821 (
            .O(N__8699),
            .I(N__8695));
    InMux I__1820 (
            .O(N__8698),
            .I(N__8692));
    Span4Mux_h I__1819 (
            .O(N__8695),
            .I(N__8689));
    LocalMux I__1818 (
            .O(N__8692),
            .I(N__8684));
    Span4Mux_v I__1817 (
            .O(N__8689),
            .I(N__8684));
    Odrv4 I__1816 (
            .O(N__8684),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ));
    InMux I__1815 (
            .O(N__8681),
            .I(N__8675));
    InMux I__1814 (
            .O(N__8680),
            .I(N__8675));
    LocalMux I__1813 (
            .O(N__8675),
            .I(\U712_REG_SM.N_95 ));
    IoInMux I__1812 (
            .O(N__8672),
            .I(N__8669));
    LocalMux I__1811 (
            .O(N__8669),
            .I(N__8666));
    Span4Mux_s3_v I__1810 (
            .O(N__8666),
            .I(N__8663));
    Span4Mux_v I__1809 (
            .O(N__8663),
            .I(N__8660));
    Span4Mux_v I__1808 (
            .O(N__8660),
            .I(N__8656));
    CascadeMux I__1807 (
            .O(N__8659),
            .I(N__8653));
    Sp12to4 I__1806 (
            .O(N__8656),
            .I(N__8650));
    InMux I__1805 (
            .O(N__8653),
            .I(N__8647));
    Odrv12 I__1804 (
            .O(N__8650),
            .I(UDSn_c));
    LocalMux I__1803 (
            .O(N__8647),
            .I(UDSn_c));
    InMux I__1802 (
            .O(N__8642),
            .I(N__8639));
    LocalMux I__1801 (
            .O(N__8639),
            .I(\U712_REG_SM.N_433 ));
    IoInMux I__1800 (
            .O(N__8636),
            .I(N__8633));
    LocalMux I__1799 (
            .O(N__8633),
            .I(N__8630));
    Odrv12 I__1798 (
            .O(N__8630),
            .I(RESETn_c_i));
    CascadeMux I__1797 (
            .O(N__8627),
            .I(N__8624));
    InMux I__1796 (
            .O(N__8624),
            .I(N__8621));
    LocalMux I__1795 (
            .O(N__8621),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ));
    IoInMux I__1794 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__1793 (
            .O(N__8615),
            .I(N__8612));
    Span12Mux_s3_h I__1792 (
            .O(N__8612),
            .I(N__8609));
    Span12Mux_h I__1791 (
            .O(N__8609),
            .I(N__8606));
    Odrv12 I__1790 (
            .O(N__8606),
            .I(CMA_c_3));
    InMux I__1789 (
            .O(N__8603),
            .I(N__8600));
    LocalMux I__1788 (
            .O(N__8600),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ));
    IoInMux I__1787 (
            .O(N__8597),
            .I(N__8594));
    LocalMux I__1786 (
            .O(N__8594),
            .I(N__8591));
    Span12Mux_s3_h I__1785 (
            .O(N__8591),
            .I(N__8588));
    Span12Mux_h I__1784 (
            .O(N__8588),
            .I(N__8585));
    Odrv12 I__1783 (
            .O(N__8585),
            .I(CMA_c_4));
    InMux I__1782 (
            .O(N__8582),
            .I(N__8577));
    InMux I__1781 (
            .O(N__8581),
            .I(N__8572));
    InMux I__1780 (
            .O(N__8580),
            .I(N__8572));
    LocalMux I__1779 (
            .O(N__8577),
            .I(N__8564));
    LocalMux I__1778 (
            .O(N__8572),
            .I(N__8564));
    InMux I__1777 (
            .O(N__8571),
            .I(N__8557));
    InMux I__1776 (
            .O(N__8570),
            .I(N__8557));
    InMux I__1775 (
            .O(N__8569),
            .I(N__8557));
    Span4Mux_h I__1774 (
            .O(N__8564),
            .I(N__8552));
    LocalMux I__1773 (
            .O(N__8557),
            .I(N__8552));
    Span4Mux_h I__1772 (
            .O(N__8552),
            .I(N__8545));
    InMux I__1771 (
            .O(N__8551),
            .I(N__8542));
    InMux I__1770 (
            .O(N__8550),
            .I(N__8539));
    InMux I__1769 (
            .O(N__8549),
            .I(N__8536));
    InMux I__1768 (
            .O(N__8548),
            .I(N__8533));
    Odrv4 I__1767 (
            .O(N__8545),
            .I(\U712_CHIP_RAM.N_297 ));
    LocalMux I__1766 (
            .O(N__8542),
            .I(\U712_CHIP_RAM.N_297 ));
    LocalMux I__1765 (
            .O(N__8539),
            .I(\U712_CHIP_RAM.N_297 ));
    LocalMux I__1764 (
            .O(N__8536),
            .I(\U712_CHIP_RAM.N_297 ));
    LocalMux I__1763 (
            .O(N__8533),
            .I(\U712_CHIP_RAM.N_297 ));
    CascadeMux I__1762 (
            .O(N__8522),
            .I(N__8516));
    CascadeMux I__1761 (
            .O(N__8521),
            .I(N__8513));
    CascadeMux I__1760 (
            .O(N__8520),
            .I(N__8508));
    CascadeMux I__1759 (
            .O(N__8519),
            .I(N__8505));
    InMux I__1758 (
            .O(N__8516),
            .I(N__8501));
    InMux I__1757 (
            .O(N__8513),
            .I(N__8498));
    InMux I__1756 (
            .O(N__8512),
            .I(N__8493));
    InMux I__1755 (
            .O(N__8511),
            .I(N__8493));
    InMux I__1754 (
            .O(N__8508),
            .I(N__8490));
    InMux I__1753 (
            .O(N__8505),
            .I(N__8485));
    InMux I__1752 (
            .O(N__8504),
            .I(N__8485));
    LocalMux I__1751 (
            .O(N__8501),
            .I(N__8480));
    LocalMux I__1750 (
            .O(N__8498),
            .I(N__8480));
    LocalMux I__1749 (
            .O(N__8493),
            .I(N__8473));
    LocalMux I__1748 (
            .O(N__8490),
            .I(N__8473));
    LocalMux I__1747 (
            .O(N__8485),
            .I(N__8473));
    Span4Mux_h I__1746 (
            .O(N__8480),
            .I(N__8470));
    Odrv4 I__1745 (
            .O(N__8473),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    Odrv4 I__1744 (
            .O(N__8470),
            .I(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ));
    InMux I__1743 (
            .O(N__8465),
            .I(N__8462));
    LocalMux I__1742 (
            .O(N__8462),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ));
    IoInMux I__1741 (
            .O(N__8459),
            .I(N__8456));
    LocalMux I__1740 (
            .O(N__8456),
            .I(N__8453));
    IoSpan4Mux I__1739 (
            .O(N__8453),
            .I(N__8450));
    Span4Mux_s1_h I__1738 (
            .O(N__8450),
            .I(N__8447));
    Sp12to4 I__1737 (
            .O(N__8447),
            .I(N__8444));
    Span12Mux_h I__1736 (
            .O(N__8444),
            .I(N__8441));
    Odrv12 I__1735 (
            .O(N__8441),
            .I(CMA_c_6));
    InMux I__1734 (
            .O(N__8438),
            .I(N__8435));
    LocalMux I__1733 (
            .O(N__8435),
            .I(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ));
    InMux I__1732 (
            .O(N__8432),
            .I(N__8429));
    LocalMux I__1731 (
            .O(N__8429),
            .I(N__8426));
    Odrv4 I__1730 (
            .O(N__8426),
            .I(\U712_CHIP_RAM.DMA_AZ0Z1 ));
    InMux I__1729 (
            .O(N__8423),
            .I(N__8420));
    LocalMux I__1728 (
            .O(N__8420),
            .I(N__8417));
    Span4Mux_v I__1727 (
            .O(N__8417),
            .I(N__8414));
    Odrv4 I__1726 (
            .O(N__8414),
            .I(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ));
    InMux I__1725 (
            .O(N__8411),
            .I(N__8408));
    LocalMux I__1724 (
            .O(N__8408),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ));
    InMux I__1723 (
            .O(N__8405),
            .I(N__8402));
    LocalMux I__1722 (
            .O(N__8402),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ));
    InMux I__1721 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__1720 (
            .O(N__8396),
            .I(\U712_BYTE_ENABLE.N_451 ));
    IoInMux I__1719 (
            .O(N__8393),
            .I(N__8390));
    LocalMux I__1718 (
            .O(N__8390),
            .I(N__8387));
    Span4Mux_s3_v I__1717 (
            .O(N__8387),
            .I(N__8384));
    Span4Mux_h I__1716 (
            .O(N__8384),
            .I(N__8381));
    Sp12to4 I__1715 (
            .O(N__8381),
            .I(N__8378));
    Span12Mux_s10_v I__1714 (
            .O(N__8378),
            .I(N__8375));
    Odrv12 I__1713 (
            .O(N__8375),
            .I(N_211_i));
    CascadeMux I__1712 (
            .O(N__8372),
            .I(\U712_BYTE_ENABLE.N_410_cascade_ ));
    IoInMux I__1711 (
            .O(N__8369),
            .I(N__8366));
    LocalMux I__1710 (
            .O(N__8366),
            .I(N__8363));
    Span12Mux_s4_h I__1709 (
            .O(N__8363),
            .I(N__8360));
    Span12Mux_h I__1708 (
            .O(N__8360),
            .I(N__8357));
    Span12Mux_v I__1707 (
            .O(N__8357),
            .I(N__8354));
    Odrv12 I__1706 (
            .O(N__8354),
            .I(N_148_i));
    InMux I__1705 (
            .O(N__8351),
            .I(N__8345));
    InMux I__1704 (
            .O(N__8350),
            .I(N__8345));
    LocalMux I__1703 (
            .O(N__8345),
            .I(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0 ));
    InMux I__1702 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__1701 (
            .O(N__8339),
            .I(N__8333));
    InMux I__1700 (
            .O(N__8338),
            .I(N__8330));
    InMux I__1699 (
            .O(N__8337),
            .I(N__8326));
    InMux I__1698 (
            .O(N__8336),
            .I(N__8323));
    Span4Mux_h I__1697 (
            .O(N__8333),
            .I(N__8320));
    LocalMux I__1696 (
            .O(N__8330),
            .I(N__8317));
    InMux I__1695 (
            .O(N__8329),
            .I(N__8314));
    LocalMux I__1694 (
            .O(N__8326),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1693 (
            .O(N__8323),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__1692 (
            .O(N__8320),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    Odrv4 I__1691 (
            .O(N__8317),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    LocalMux I__1690 (
            .O(N__8314),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_1 ));
    InMux I__1689 (
            .O(N__8303),
            .I(N__8300));
    LocalMux I__1688 (
            .O(N__8300),
            .I(N__8291));
    InMux I__1687 (
            .O(N__8299),
            .I(N__8288));
    CascadeMux I__1686 (
            .O(N__8298),
            .I(N__8285));
    CascadeMux I__1685 (
            .O(N__8297),
            .I(N__8281));
    CascadeMux I__1684 (
            .O(N__8296),
            .I(N__8277));
    InMux I__1683 (
            .O(N__8295),
            .I(N__8270));
    InMux I__1682 (
            .O(N__8294),
            .I(N__8270));
    Span4Mux_h I__1681 (
            .O(N__8291),
            .I(N__8267));
    LocalMux I__1680 (
            .O(N__8288),
            .I(N__8264));
    InMux I__1679 (
            .O(N__8285),
            .I(N__8261));
    InMux I__1678 (
            .O(N__8284),
            .I(N__8258));
    InMux I__1677 (
            .O(N__8281),
            .I(N__8253));
    InMux I__1676 (
            .O(N__8280),
            .I(N__8253));
    InMux I__1675 (
            .O(N__8277),
            .I(N__8250));
    InMux I__1674 (
            .O(N__8276),
            .I(N__8245));
    InMux I__1673 (
            .O(N__8275),
            .I(N__8245));
    LocalMux I__1672 (
            .O(N__8270),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1671 (
            .O(N__8267),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    Odrv4 I__1670 (
            .O(N__8264),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1669 (
            .O(N__8261),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1668 (
            .O(N__8258),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1667 (
            .O(N__8253),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1666 (
            .O(N__8250),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    LocalMux I__1665 (
            .O(N__8245),
            .I(\U712_REG_SM.C3_SYNCZ0Z_1 ));
    InMux I__1664 (
            .O(N__8228),
            .I(N__8222));
    CascadeMux I__1663 (
            .O(N__8227),
            .I(N__8217));
    CascadeMux I__1662 (
            .O(N__8226),
            .I(N__8214));
    InMux I__1661 (
            .O(N__8225),
            .I(N__8210));
    LocalMux I__1660 (
            .O(N__8222),
            .I(N__8207));
    InMux I__1659 (
            .O(N__8221),
            .I(N__8202));
    InMux I__1658 (
            .O(N__8220),
            .I(N__8202));
    InMux I__1657 (
            .O(N__8217),
            .I(N__8197));
    InMux I__1656 (
            .O(N__8214),
            .I(N__8197));
    InMux I__1655 (
            .O(N__8213),
            .I(N__8194));
    LocalMux I__1654 (
            .O(N__8210),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    Odrv4 I__1653 (
            .O(N__8207),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1652 (
            .O(N__8202),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1651 (
            .O(N__8197),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    LocalMux I__1650 (
            .O(N__8194),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_8 ));
    CascadeMux I__1649 (
            .O(N__8183),
            .I(\U712_REG_SM.N_95_cascade_ ));
    InMux I__1648 (
            .O(N__8180),
            .I(N__8177));
    LocalMux I__1647 (
            .O(N__8177),
            .I(\U712_REG_SM.N_432 ));
    IoInMux I__1646 (
            .O(N__8174),
            .I(N__8171));
    LocalMux I__1645 (
            .O(N__8171),
            .I(N__8168));
    Span12Mux_s0_v I__1644 (
            .O(N__8168),
            .I(N__8165));
    Span12Mux_h I__1643 (
            .O(N__8165),
            .I(N__8161));
    InMux I__1642 (
            .O(N__8164),
            .I(N__8158));
    Odrv12 I__1641 (
            .O(N__8161),
            .I(LDSn_c));
    LocalMux I__1640 (
            .O(N__8158),
            .I(LDSn_c));
    CascadeMux I__1639 (
            .O(N__8153),
            .I(N__8146));
    CascadeMux I__1638 (
            .O(N__8152),
            .I(N__8143));
    CascadeMux I__1637 (
            .O(N__8151),
            .I(N__8140));
    InMux I__1636 (
            .O(N__8150),
            .I(N__8134));
    InMux I__1635 (
            .O(N__8149),
            .I(N__8134));
    InMux I__1634 (
            .O(N__8146),
            .I(N__8131));
    InMux I__1633 (
            .O(N__8143),
            .I(N__8126));
    InMux I__1632 (
            .O(N__8140),
            .I(N__8126));
    InMux I__1631 (
            .O(N__8139),
            .I(N__8121));
    LocalMux I__1630 (
            .O(N__8134),
            .I(N__8106));
    LocalMux I__1629 (
            .O(N__8131),
            .I(N__8106));
    LocalMux I__1628 (
            .O(N__8126),
            .I(N__8106));
    InMux I__1627 (
            .O(N__8125),
            .I(N__8101));
    InMux I__1626 (
            .O(N__8124),
            .I(N__8101));
    LocalMux I__1625 (
            .O(N__8121),
            .I(N__8098));
    InMux I__1624 (
            .O(N__8120),
            .I(N__8095));
    InMux I__1623 (
            .O(N__8119),
            .I(N__8092));
    InMux I__1622 (
            .O(N__8118),
            .I(N__8089));
    InMux I__1621 (
            .O(N__8117),
            .I(N__8082));
    InMux I__1620 (
            .O(N__8116),
            .I(N__8082));
    InMux I__1619 (
            .O(N__8115),
            .I(N__8082));
    InMux I__1618 (
            .O(N__8114),
            .I(N__8077));
    InMux I__1617 (
            .O(N__8113),
            .I(N__8077));
    Span4Mux_v I__1616 (
            .O(N__8106),
            .I(N__8074));
    LocalMux I__1615 (
            .O(N__8101),
            .I(N__8071));
    Odrv12 I__1614 (
            .O(N__8098),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1613 (
            .O(N__8095),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1612 (
            .O(N__8092),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1611 (
            .O(N__8089),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1610 (
            .O(N__8082),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    LocalMux I__1609 (
            .O(N__8077),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1608 (
            .O(N__8074),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    Odrv4 I__1607 (
            .O(N__8071),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ));
    InMux I__1606 (
            .O(N__8054),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ));
    CascadeMux I__1605 (
            .O(N__8051),
            .I(N__8047));
    CascadeMux I__1604 (
            .O(N__8050),
            .I(N__8044));
    InMux I__1603 (
            .O(N__8047),
            .I(N__8035));
    InMux I__1602 (
            .O(N__8044),
            .I(N__8031));
    InMux I__1601 (
            .O(N__8043),
            .I(N__8026));
    InMux I__1600 (
            .O(N__8042),
            .I(N__8026));
    InMux I__1599 (
            .O(N__8041),
            .I(N__8023));
    InMux I__1598 (
            .O(N__8040),
            .I(N__8017));
    InMux I__1597 (
            .O(N__8039),
            .I(N__8011));
    InMux I__1596 (
            .O(N__8038),
            .I(N__8011));
    LocalMux I__1595 (
            .O(N__8035),
            .I(N__8008));
    CascadeMux I__1594 (
            .O(N__8034),
            .I(N__8001));
    LocalMux I__1593 (
            .O(N__8031),
            .I(N__7997));
    LocalMux I__1592 (
            .O(N__8026),
            .I(N__7992));
    LocalMux I__1591 (
            .O(N__8023),
            .I(N__7992));
    InMux I__1590 (
            .O(N__8022),
            .I(N__7985));
    InMux I__1589 (
            .O(N__8021),
            .I(N__7985));
    InMux I__1588 (
            .O(N__8020),
            .I(N__7985));
    LocalMux I__1587 (
            .O(N__8017),
            .I(N__7977));
    InMux I__1586 (
            .O(N__8016),
            .I(N__7974));
    LocalMux I__1585 (
            .O(N__8011),
            .I(N__7969));
    Span4Mux_v I__1584 (
            .O(N__8008),
            .I(N__7969));
    InMux I__1583 (
            .O(N__8007),
            .I(N__7960));
    InMux I__1582 (
            .O(N__8006),
            .I(N__7960));
    InMux I__1581 (
            .O(N__8005),
            .I(N__7960));
    InMux I__1580 (
            .O(N__8004),
            .I(N__7960));
    InMux I__1579 (
            .O(N__8001),
            .I(N__7955));
    InMux I__1578 (
            .O(N__8000),
            .I(N__7955));
    Span4Mux_h I__1577 (
            .O(N__7997),
            .I(N__7948));
    Span4Mux_v I__1576 (
            .O(N__7992),
            .I(N__7948));
    LocalMux I__1575 (
            .O(N__7985),
            .I(N__7948));
    InMux I__1574 (
            .O(N__7984),
            .I(N__7941));
    InMux I__1573 (
            .O(N__7983),
            .I(N__7941));
    InMux I__1572 (
            .O(N__7982),
            .I(N__7941));
    InMux I__1571 (
            .O(N__7981),
            .I(N__7936));
    InMux I__1570 (
            .O(N__7980),
            .I(N__7936));
    Odrv4 I__1569 (
            .O(N__7977),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1568 (
            .O(N__7974),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1567 (
            .O(N__7969),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1566 (
            .O(N__7960),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1565 (
            .O(N__7955),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    Odrv4 I__1564 (
            .O(N__7948),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1563 (
            .O(N__7941),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    LocalMux I__1562 (
            .O(N__7936),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ));
    CascadeMux I__1561 (
            .O(N__7919),
            .I(N__7916));
    InMux I__1560 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__1559 (
            .O(N__7913),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ));
    InMux I__1558 (
            .O(N__7910),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ));
    CascadeMux I__1557 (
            .O(N__7907),
            .I(N__7902));
    InMux I__1556 (
            .O(N__7906),
            .I(N__7898));
    CascadeMux I__1555 (
            .O(N__7905),
            .I(N__7894));
    InMux I__1554 (
            .O(N__7902),
            .I(N__7889));
    InMux I__1553 (
            .O(N__7901),
            .I(N__7889));
    LocalMux I__1552 (
            .O(N__7898),
            .I(N__7885));
    InMux I__1551 (
            .O(N__7897),
            .I(N__7880));
    InMux I__1550 (
            .O(N__7894),
            .I(N__7880));
    LocalMux I__1549 (
            .O(N__7889),
            .I(N__7877));
    InMux I__1548 (
            .O(N__7888),
            .I(N__7869));
    Span4Mux_h I__1547 (
            .O(N__7885),
            .I(N__7866));
    LocalMux I__1546 (
            .O(N__7880),
            .I(N__7863));
    Span4Mux_h I__1545 (
            .O(N__7877),
            .I(N__7860));
    InMux I__1544 (
            .O(N__7876),
            .I(N__7853));
    InMux I__1543 (
            .O(N__7875),
            .I(N__7853));
    InMux I__1542 (
            .O(N__7874),
            .I(N__7853));
    InMux I__1541 (
            .O(N__7873),
            .I(N__7848));
    InMux I__1540 (
            .O(N__7872),
            .I(N__7848));
    LocalMux I__1539 (
            .O(N__7869),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1538 (
            .O(N__7866),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1537 (
            .O(N__7863),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    Odrv4 I__1536 (
            .O(N__7860),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1535 (
            .O(N__7853),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    LocalMux I__1534 (
            .O(N__7848),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ));
    InMux I__1533 (
            .O(N__7835),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ));
    InMux I__1532 (
            .O(N__7832),
            .I(N__7828));
    InMux I__1531 (
            .O(N__7831),
            .I(N__7825));
    LocalMux I__1530 (
            .O(N__7828),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    LocalMux I__1529 (
            .O(N__7825),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ));
    InMux I__1528 (
            .O(N__7820),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ));
    InMux I__1527 (
            .O(N__7817),
            .I(N__7813));
    InMux I__1526 (
            .O(N__7816),
            .I(N__7810));
    LocalMux I__1525 (
            .O(N__7813),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    LocalMux I__1524 (
            .O(N__7810),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ));
    InMux I__1523 (
            .O(N__7805),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ));
    InMux I__1522 (
            .O(N__7802),
            .I(N__7798));
    InMux I__1521 (
            .O(N__7801),
            .I(N__7795));
    LocalMux I__1520 (
            .O(N__7798),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    LocalMux I__1519 (
            .O(N__7795),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ));
    InMux I__1518 (
            .O(N__7790),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ));
    InMux I__1517 (
            .O(N__7787),
            .I(N__7772));
    InMux I__1516 (
            .O(N__7786),
            .I(N__7772));
    InMux I__1515 (
            .O(N__7785),
            .I(N__7772));
    InMux I__1514 (
            .O(N__7784),
            .I(N__7772));
    InMux I__1513 (
            .O(N__7783),
            .I(N__7769));
    InMux I__1512 (
            .O(N__7782),
            .I(N__7764));
    InMux I__1511 (
            .O(N__7781),
            .I(N__7764));
    LocalMux I__1510 (
            .O(N__7772),
            .I(\U712_CHIP_RAM.N_200 ));
    LocalMux I__1509 (
            .O(N__7769),
            .I(\U712_CHIP_RAM.N_200 ));
    LocalMux I__1508 (
            .O(N__7764),
            .I(\U712_CHIP_RAM.N_200 ));
    InMux I__1507 (
            .O(N__7757),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ));
    CascadeMux I__1506 (
            .O(N__7754),
            .I(N__7750));
    InMux I__1505 (
            .O(N__7753),
            .I(N__7747));
    InMux I__1504 (
            .O(N__7750),
            .I(N__7744));
    LocalMux I__1503 (
            .O(N__7747),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    LocalMux I__1502 (
            .O(N__7744),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ));
    CEMux I__1501 (
            .O(N__7739),
            .I(N__7736));
    LocalMux I__1500 (
            .O(N__7736),
            .I(N__7733));
    Span4Mux_v I__1499 (
            .O(N__7733),
            .I(N__7729));
    CEMux I__1498 (
            .O(N__7732),
            .I(N__7726));
    Span4Mux_v I__1497 (
            .O(N__7729),
            .I(N__7721));
    LocalMux I__1496 (
            .O(N__7726),
            .I(N__7721));
    Span4Mux_h I__1495 (
            .O(N__7721),
            .I(N__7718));
    Odrv4 I__1494 (
            .O(N__7718),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ));
    InMux I__1493 (
            .O(N__7715),
            .I(N__7712));
    LocalMux I__1492 (
            .O(N__7712),
            .I(N__7709));
    Odrv12 I__1491 (
            .O(N__7709),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ));
    CascadeMux I__1490 (
            .O(N__7706),
            .I(\U712_CHIP_RAM.N_294_cascade_ ));
    CascadeMux I__1489 (
            .O(N__7703),
            .I(N__7700));
    InMux I__1488 (
            .O(N__7700),
            .I(N__7696));
    InMux I__1487 (
            .O(N__7699),
            .I(N__7693));
    LocalMux I__1486 (
            .O(N__7696),
            .I(N__7687));
    LocalMux I__1485 (
            .O(N__7693),
            .I(N__7687));
    InMux I__1484 (
            .O(N__7692),
            .I(N__7679));
    Span4Mux_h I__1483 (
            .O(N__7687),
            .I(N__7672));
    InMux I__1482 (
            .O(N__7686),
            .I(N__7669));
    InMux I__1481 (
            .O(N__7685),
            .I(N__7664));
    InMux I__1480 (
            .O(N__7684),
            .I(N__7664));
    InMux I__1479 (
            .O(N__7683),
            .I(N__7659));
    InMux I__1478 (
            .O(N__7682),
            .I(N__7659));
    LocalMux I__1477 (
            .O(N__7679),
            .I(N__7656));
    InMux I__1476 (
            .O(N__7678),
            .I(N__7651));
    InMux I__1475 (
            .O(N__7677),
            .I(N__7651));
    InMux I__1474 (
            .O(N__7676),
            .I(N__7646));
    InMux I__1473 (
            .O(N__7675),
            .I(N__7646));
    Odrv4 I__1472 (
            .O(N__7672),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__1471 (
            .O(N__7669),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__1470 (
            .O(N__7664),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__1469 (
            .O(N__7659),
            .I(\U712_CHIP_RAM.N_288 ));
    Odrv4 I__1468 (
            .O(N__7656),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__1467 (
            .O(N__7651),
            .I(\U712_CHIP_RAM.N_288 ));
    LocalMux I__1466 (
            .O(N__7646),
            .I(\U712_CHIP_RAM.N_288 ));
    CascadeMux I__1465 (
            .O(N__7631),
            .I(\U712_CHIP_RAM.N_469_cascade_ ));
    InMux I__1464 (
            .O(N__7628),
            .I(N__7624));
    InMux I__1463 (
            .O(N__7627),
            .I(N__7619));
    LocalMux I__1462 (
            .O(N__7624),
            .I(N__7616));
    InMux I__1461 (
            .O(N__7623),
            .I(N__7613));
    InMux I__1460 (
            .O(N__7622),
            .I(N__7610));
    LocalMux I__1459 (
            .O(N__7619),
            .I(\U712_CHIP_RAM.N_557 ));
    Odrv4 I__1458 (
            .O(N__7616),
            .I(\U712_CHIP_RAM.N_557 ));
    LocalMux I__1457 (
            .O(N__7613),
            .I(\U712_CHIP_RAM.N_557 ));
    LocalMux I__1456 (
            .O(N__7610),
            .I(\U712_CHIP_RAM.N_557 ));
    InMux I__1455 (
            .O(N__7601),
            .I(N__7593));
    InMux I__1454 (
            .O(N__7600),
            .I(N__7593));
    InMux I__1453 (
            .O(N__7599),
            .I(N__7582));
    InMux I__1452 (
            .O(N__7598),
            .I(N__7582));
    LocalMux I__1451 (
            .O(N__7593),
            .I(N__7577));
    CascadeMux I__1450 (
            .O(N__7592),
            .I(N__7571));
    InMux I__1449 (
            .O(N__7591),
            .I(N__7564));
    InMux I__1448 (
            .O(N__7590),
            .I(N__7564));
    InMux I__1447 (
            .O(N__7589),
            .I(N__7559));
    InMux I__1446 (
            .O(N__7588),
            .I(N__7559));
    InMux I__1445 (
            .O(N__7587),
            .I(N__7556));
    LocalMux I__1444 (
            .O(N__7582),
            .I(N__7553));
    InMux I__1443 (
            .O(N__7581),
            .I(N__7548));
    InMux I__1442 (
            .O(N__7580),
            .I(N__7548));
    Span4Mux_h I__1441 (
            .O(N__7577),
            .I(N__7545));
    InMux I__1440 (
            .O(N__7576),
            .I(N__7538));
    InMux I__1439 (
            .O(N__7575),
            .I(N__7538));
    InMux I__1438 (
            .O(N__7574),
            .I(N__7538));
    InMux I__1437 (
            .O(N__7571),
            .I(N__7531));
    InMux I__1436 (
            .O(N__7570),
            .I(N__7531));
    InMux I__1435 (
            .O(N__7569),
            .I(N__7531));
    LocalMux I__1434 (
            .O(N__7564),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1433 (
            .O(N__7559),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1432 (
            .O(N__7556),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1431 (
            .O(N__7553),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1430 (
            .O(N__7548),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    Odrv4 I__1429 (
            .O(N__7545),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1428 (
            .O(N__7538),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    LocalMux I__1427 (
            .O(N__7531),
            .I(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ));
    InMux I__1426 (
            .O(N__7514),
            .I(N__7511));
    LocalMux I__1425 (
            .O(N__7511),
            .I(\U712_CHIP_RAM.N_555 ));
    CascadeMux I__1424 (
            .O(N__7508),
            .I(\U712_CHIP_RAM.N_309_cascade_ ));
    InMux I__1423 (
            .O(N__7505),
            .I(N__7502));
    LocalMux I__1422 (
            .O(N__7502),
            .I(\U712_CHIP_RAM.N_387 ));
    CascadeMux I__1421 (
            .O(N__7499),
            .I(\U712_CHIP_RAM.N_200_cascade_ ));
    InMux I__1420 (
            .O(N__7496),
            .I(N__7493));
    LocalMux I__1419 (
            .O(N__7493),
            .I(\U712_CHIP_RAM.N_309 ));
    InMux I__1418 (
            .O(N__7490),
            .I(N__7486));
    CascadeMux I__1417 (
            .O(N__7489),
            .I(N__7482));
    LocalMux I__1416 (
            .O(N__7486),
            .I(N__7479));
    InMux I__1415 (
            .O(N__7485),
            .I(N__7474));
    InMux I__1414 (
            .O(N__7482),
            .I(N__7474));
    Odrv4 I__1413 (
            .O(N__7479),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    LocalMux I__1412 (
            .O(N__7474),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ));
    InMux I__1411 (
            .O(N__7469),
            .I(N__7463));
    InMux I__1410 (
            .O(N__7468),
            .I(N__7460));
    InMux I__1409 (
            .O(N__7467),
            .I(N__7457));
    InMux I__1408 (
            .O(N__7466),
            .I(N__7454));
    LocalMux I__1407 (
            .O(N__7463),
            .I(N__7451));
    LocalMux I__1406 (
            .O(N__7460),
            .I(N__7448));
    LocalMux I__1405 (
            .O(N__7457),
            .I(N__7443));
    LocalMux I__1404 (
            .O(N__7454),
            .I(N__7443));
    Span4Mux_h I__1403 (
            .O(N__7451),
            .I(N__7439));
    Span4Mux_h I__1402 (
            .O(N__7448),
            .I(N__7436));
    Span4Mux_v I__1401 (
            .O(N__7443),
            .I(N__7433));
    InMux I__1400 (
            .O(N__7442),
            .I(N__7430));
    Odrv4 I__1399 (
            .O(N__7439),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1398 (
            .O(N__7436),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    Odrv4 I__1397 (
            .O(N__7433),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    LocalMux I__1396 (
            .O(N__7430),
            .I(\U712_CHIP_RAM.WRITE_CYCLEZ0 ));
    InMux I__1395 (
            .O(N__7421),
            .I(N__7416));
    InMux I__1394 (
            .O(N__7420),
            .I(N__7413));
    InMux I__1393 (
            .O(N__7419),
            .I(N__7410));
    LocalMux I__1392 (
            .O(N__7416),
            .I(N__7407));
    LocalMux I__1391 (
            .O(N__7413),
            .I(N__7404));
    LocalMux I__1390 (
            .O(N__7410),
            .I(N__7401));
    Span4Mux_h I__1389 (
            .O(N__7407),
            .I(N__7398));
    Span4Mux_h I__1388 (
            .O(N__7404),
            .I(N__7395));
    Odrv4 I__1387 (
            .O(N__7401),
            .I(\U712_CHIP_RAM.N_285 ));
    Odrv4 I__1386 (
            .O(N__7398),
            .I(\U712_CHIP_RAM.N_285 ));
    Odrv4 I__1385 (
            .O(N__7395),
            .I(\U712_CHIP_RAM.N_285 ));
    CascadeMux I__1384 (
            .O(N__7388),
            .I(\U712_CHIP_RAM.N_285_cascade_ ));
    InMux I__1383 (
            .O(N__7385),
            .I(N__7382));
    LocalMux I__1382 (
            .O(N__7382),
            .I(N__7379));
    Span4Mux_h I__1381 (
            .O(N__7379),
            .I(N__7371));
    InMux I__1380 (
            .O(N__7378),
            .I(N__7366));
    InMux I__1379 (
            .O(N__7377),
            .I(N__7366));
    InMux I__1378 (
            .O(N__7376),
            .I(N__7363));
    InMux I__1377 (
            .O(N__7375),
            .I(N__7358));
    InMux I__1376 (
            .O(N__7374),
            .I(N__7358));
    Odrv4 I__1375 (
            .O(N__7371),
            .I(\U712_CHIP_RAM.N_293 ));
    LocalMux I__1374 (
            .O(N__7366),
            .I(\U712_CHIP_RAM.N_293 ));
    LocalMux I__1373 (
            .O(N__7363),
            .I(\U712_CHIP_RAM.N_293 ));
    LocalMux I__1372 (
            .O(N__7358),
            .I(\U712_CHIP_RAM.N_293 ));
    CascadeMux I__1371 (
            .O(N__7349),
            .I(N__7346));
    InMux I__1370 (
            .O(N__7346),
            .I(N__7343));
    LocalMux I__1369 (
            .O(N__7343),
            .I(N__7340));
    Span4Mux_h I__1368 (
            .O(N__7340),
            .I(N__7337));
    Odrv4 I__1367 (
            .O(N__7337),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2 ));
    CascadeMux I__1366 (
            .O(N__7334),
            .I(N__7330));
    CascadeMux I__1365 (
            .O(N__7333),
            .I(N__7325));
    InMux I__1364 (
            .O(N__7330),
            .I(N__7320));
    InMux I__1363 (
            .O(N__7329),
            .I(N__7317));
    InMux I__1362 (
            .O(N__7328),
            .I(N__7314));
    InMux I__1361 (
            .O(N__7325),
            .I(N__7309));
    InMux I__1360 (
            .O(N__7324),
            .I(N__7309));
    InMux I__1359 (
            .O(N__7323),
            .I(N__7304));
    LocalMux I__1358 (
            .O(N__7320),
            .I(N__7299));
    LocalMux I__1357 (
            .O(N__7317),
            .I(N__7299));
    LocalMux I__1356 (
            .O(N__7314),
            .I(N__7294));
    LocalMux I__1355 (
            .O(N__7309),
            .I(N__7294));
    CascadeMux I__1354 (
            .O(N__7308),
            .I(N__7287));
    InMux I__1353 (
            .O(N__7307),
            .I(N__7282));
    LocalMux I__1352 (
            .O(N__7304),
            .I(N__7277));
    Span4Mux_v I__1351 (
            .O(N__7299),
            .I(N__7277));
    Span4Mux_v I__1350 (
            .O(N__7294),
            .I(N__7274));
    InMux I__1349 (
            .O(N__7293),
            .I(N__7265));
    InMux I__1348 (
            .O(N__7292),
            .I(N__7265));
    InMux I__1347 (
            .O(N__7291),
            .I(N__7265));
    InMux I__1346 (
            .O(N__7290),
            .I(N__7265));
    InMux I__1345 (
            .O(N__7287),
            .I(N__7258));
    InMux I__1344 (
            .O(N__7286),
            .I(N__7258));
    InMux I__1343 (
            .O(N__7285),
            .I(N__7258));
    LocalMux I__1342 (
            .O(N__7282),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1341 (
            .O(N__7277),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    Odrv4 I__1340 (
            .O(N__7274),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1339 (
            .O(N__7265),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    LocalMux I__1338 (
            .O(N__7258),
            .I(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ));
    InMux I__1337 (
            .O(N__7247),
            .I(N__7244));
    LocalMux I__1336 (
            .O(N__7244),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ));
    InMux I__1335 (
            .O(N__7241),
            .I(bfn_12_9_0_));
    InMux I__1334 (
            .O(N__7238),
            .I(N__7235));
    LocalMux I__1333 (
            .O(N__7235),
            .I(N__7232));
    Span4Mux_v I__1332 (
            .O(N__7232),
            .I(N__7229));
    Span4Mux_h I__1331 (
            .O(N__7229),
            .I(N__7226));
    Sp12to4 I__1330 (
            .O(N__7226),
            .I(N__7223));
    Span12Mux_h I__1329 (
            .O(N__7223),
            .I(N__7220));
    Span12Mux_v I__1328 (
            .O(N__7220),
            .I(N__7217));
    Odrv12 I__1327 (
            .O(N__7217),
            .I(A_c_3));
    InMux I__1326 (
            .O(N__7214),
            .I(N__7211));
    LocalMux I__1325 (
            .O(N__7211),
            .I(N__7208));
    Span4Mux_h I__1324 (
            .O(N__7208),
            .I(N__7205));
    Odrv4 I__1323 (
            .O(N__7205),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ));
    InMux I__1322 (
            .O(N__7202),
            .I(N__7199));
    LocalMux I__1321 (
            .O(N__7199),
            .I(N__7196));
    Span4Mux_h I__1320 (
            .O(N__7196),
            .I(N__7193));
    Sp12to4 I__1319 (
            .O(N__7193),
            .I(N__7190));
    Span12Mux_v I__1318 (
            .O(N__7190),
            .I(N__7187));
    Span12Mux_h I__1317 (
            .O(N__7187),
            .I(N__7184));
    Odrv12 I__1316 (
            .O(N__7184),
            .I(A_c_4));
    InMux I__1315 (
            .O(N__7181),
            .I(N__7178));
    LocalMux I__1314 (
            .O(N__7178),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ));
    InMux I__1313 (
            .O(N__7175),
            .I(N__7172));
    LocalMux I__1312 (
            .O(N__7172),
            .I(N__7169));
    Span4Mux_v I__1311 (
            .O(N__7169),
            .I(N__7166));
    Span4Mux_v I__1310 (
            .O(N__7166),
            .I(N__7163));
    Sp12to4 I__1309 (
            .O(N__7163),
            .I(N__7160));
    Span12Mux_h I__1308 (
            .O(N__7160),
            .I(N__7157));
    Odrv12 I__1307 (
            .O(N__7157),
            .I(A_c_7));
    InMux I__1306 (
            .O(N__7154),
            .I(N__7151));
    LocalMux I__1305 (
            .O(N__7151),
            .I(N__7148));
    Odrv4 I__1304 (
            .O(N__7148),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ));
    InMux I__1303 (
            .O(N__7145),
            .I(N__7142));
    LocalMux I__1302 (
            .O(N__7142),
            .I(N__7139));
    Span4Mux_v I__1301 (
            .O(N__7139),
            .I(N__7136));
    Span4Mux_v I__1300 (
            .O(N__7136),
            .I(N__7133));
    Sp12to4 I__1299 (
            .O(N__7133),
            .I(N__7130));
    Span12Mux_h I__1298 (
            .O(N__7130),
            .I(N__7127));
    Odrv12 I__1297 (
            .O(N__7127),
            .I(A_c_8));
    InMux I__1296 (
            .O(N__7124),
            .I(N__7121));
    LocalMux I__1295 (
            .O(N__7121),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ));
    InMux I__1294 (
            .O(N__7118),
            .I(N__7115));
    LocalMux I__1293 (
            .O(N__7115),
            .I(N__7112));
    Span4Mux_v I__1292 (
            .O(N__7112),
            .I(N__7109));
    Span4Mux_v I__1291 (
            .O(N__7109),
            .I(N__7106));
    Sp12to4 I__1290 (
            .O(N__7106),
            .I(N__7103));
    Span12Mux_h I__1289 (
            .O(N__7103),
            .I(N__7100));
    Odrv12 I__1288 (
            .O(N__7100),
            .I(A_c_18));
    InMux I__1287 (
            .O(N__7097),
            .I(N__7094));
    LocalMux I__1286 (
            .O(N__7094),
            .I(N__7091));
    Span4Mux_h I__1285 (
            .O(N__7091),
            .I(N__7088));
    Odrv4 I__1284 (
            .O(N__7088),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ));
    InMux I__1283 (
            .O(N__7085),
            .I(N__7082));
    LocalMux I__1282 (
            .O(N__7082),
            .I(N__7079));
    Span12Mux_v I__1281 (
            .O(N__7079),
            .I(N__7076));
    Span12Mux_h I__1280 (
            .O(N__7076),
            .I(N__7073));
    Odrv12 I__1279 (
            .O(N__7073),
            .I(A_c_5));
    InMux I__1278 (
            .O(N__7070),
            .I(N__7067));
    LocalMux I__1277 (
            .O(N__7067),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ));
    CEMux I__1276 (
            .O(N__7064),
            .I(N__7061));
    LocalMux I__1275 (
            .O(N__7061),
            .I(N__7057));
    CEMux I__1274 (
            .O(N__7060),
            .I(N__7054));
    Span4Mux_v I__1273 (
            .O(N__7057),
            .I(N__7051));
    LocalMux I__1272 (
            .O(N__7054),
            .I(N__7048));
    Span4Mux_h I__1271 (
            .O(N__7051),
            .I(N__7045));
    Odrv4 I__1270 (
            .O(N__7048),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ));
    Odrv4 I__1269 (
            .O(N__7045),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ));
    InMux I__1268 (
            .O(N__7040),
            .I(N__7037));
    LocalMux I__1267 (
            .O(N__7037),
            .I(N__7033));
    InMux I__1266 (
            .O(N__7036),
            .I(N__7029));
    Span4Mux_v I__1265 (
            .O(N__7033),
            .I(N__7026));
    InMux I__1264 (
            .O(N__7032),
            .I(N__7023));
    LocalMux I__1263 (
            .O(N__7029),
            .I(N__7020));
    Sp12to4 I__1262 (
            .O(N__7026),
            .I(N__7015));
    LocalMux I__1261 (
            .O(N__7023),
            .I(N__7015));
    Span12Mux_h I__1260 (
            .O(N__7020),
            .I(N__7012));
    Span12Mux_h I__1259 (
            .O(N__7015),
            .I(N__7009));
    Span12Mux_v I__1258 (
            .O(N__7012),
            .I(N__7006));
    Span12Mux_v I__1257 (
            .O(N__7009),
            .I(N__7003));
    Odrv12 I__1256 (
            .O(N__7006),
            .I(AWEn_c));
    Odrv12 I__1255 (
            .O(N__7003),
            .I(AWEn_c));
    InMux I__1254 (
            .O(N__6998),
            .I(N__6993));
    InMux I__1253 (
            .O(N__6997),
            .I(N__6990));
    InMux I__1252 (
            .O(N__6996),
            .I(N__6987));
    LocalMux I__1251 (
            .O(N__6993),
            .I(N__6981));
    LocalMux I__1250 (
            .O(N__6990),
            .I(N__6978));
    LocalMux I__1249 (
            .O(N__6987),
            .I(N__6975));
    InMux I__1248 (
            .O(N__6986),
            .I(N__6972));
    InMux I__1247 (
            .O(N__6985),
            .I(N__6969));
    InMux I__1246 (
            .O(N__6984),
            .I(N__6963));
    Span4Mux_h I__1245 (
            .O(N__6981),
            .I(N__6960));
    Span4Mux_v I__1244 (
            .O(N__6978),
            .I(N__6953));
    Span4Mux_v I__1243 (
            .O(N__6975),
            .I(N__6953));
    LocalMux I__1242 (
            .O(N__6972),
            .I(N__6953));
    LocalMux I__1241 (
            .O(N__6969),
            .I(N__6950));
    InMux I__1240 (
            .O(N__6968),
            .I(N__6945));
    InMux I__1239 (
            .O(N__6967),
            .I(N__6945));
    InMux I__1238 (
            .O(N__6966),
            .I(N__6942));
    LocalMux I__1237 (
            .O(N__6963),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1236 (
            .O(N__6960),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1235 (
            .O(N__6953),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    Odrv4 I__1234 (
            .O(N__6950),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1233 (
            .O(N__6945),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    LocalMux I__1232 (
            .O(N__6942),
            .I(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ));
    CEMux I__1231 (
            .O(N__6929),
            .I(N__6926));
    LocalMux I__1230 (
            .O(N__6926),
            .I(N__6923));
    Span4Mux_h I__1229 (
            .O(N__6923),
            .I(N__6920));
    Odrv4 I__1228 (
            .O(N__6920),
            .I(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ));
    IoInMux I__1227 (
            .O(N__6917),
            .I(N__6914));
    LocalMux I__1226 (
            .O(N__6914),
            .I(N__6911));
    Span4Mux_s3_v I__1225 (
            .O(N__6911),
            .I(N__6908));
    Span4Mux_h I__1224 (
            .O(N__6908),
            .I(N__6905));
    Odrv4 I__1223 (
            .O(N__6905),
            .I(CONSTANT_ONE_NET));
    InMux I__1222 (
            .O(N__6902),
            .I(N__6898));
    CascadeMux I__1221 (
            .O(N__6901),
            .I(N__6894));
    LocalMux I__1220 (
            .O(N__6898),
            .I(N__6891));
    CascadeMux I__1219 (
            .O(N__6897),
            .I(N__6886));
    InMux I__1218 (
            .O(N__6894),
            .I(N__6883));
    Span4Mux_h I__1217 (
            .O(N__6891),
            .I(N__6880));
    InMux I__1216 (
            .O(N__6890),
            .I(N__6877));
    InMux I__1215 (
            .O(N__6889),
            .I(N__6874));
    InMux I__1214 (
            .O(N__6886),
            .I(N__6871));
    LocalMux I__1213 (
            .O(N__6883),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    Odrv4 I__1212 (
            .O(N__6880),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1211 (
            .O(N__6877),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1210 (
            .O(N__6874),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    LocalMux I__1209 (
            .O(N__6871),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ));
    IoInMux I__1208 (
            .O(N__6860),
            .I(N__6857));
    LocalMux I__1207 (
            .O(N__6857),
            .I(N__6854));
    Span4Mux_s2_h I__1206 (
            .O(N__6854),
            .I(N__6851));
    Span4Mux_v I__1205 (
            .O(N__6851),
            .I(N__6848));
    Sp12to4 I__1204 (
            .O(N__6848),
            .I(N__6845));
    Span12Mux_h I__1203 (
            .O(N__6845),
            .I(N__6842));
    Odrv12 I__1202 (
            .O(N__6842),
            .I(WEn_c));
    CascadeMux I__1201 (
            .O(N__6839),
            .I(N__6836));
    InMux I__1200 (
            .O(N__6836),
            .I(N__6833));
    LocalMux I__1199 (
            .O(N__6833),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ));
    InMux I__1198 (
            .O(N__6830),
            .I(N__6827));
    LocalMux I__1197 (
            .O(N__6827),
            .I(N__6824));
    Span12Mux_h I__1196 (
            .O(N__6824),
            .I(N__6821));
    Odrv12 I__1195 (
            .O(N__6821),
            .I(A_c_13));
    CascadeMux I__1194 (
            .O(N__6818),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ));
    InMux I__1193 (
            .O(N__6815),
            .I(N__6812));
    LocalMux I__1192 (
            .O(N__6812),
            .I(N__6809));
    Span12Mux_v I__1191 (
            .O(N__6809),
            .I(N__6806));
    Span12Mux_h I__1190 (
            .O(N__6806),
            .I(N__6803));
    Odrv12 I__1189 (
            .O(N__6803),
            .I(A_c_15));
    CascadeMux I__1188 (
            .O(N__6800),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ));
    InMux I__1187 (
            .O(N__6797),
            .I(N__6794));
    LocalMux I__1186 (
            .O(N__6794),
            .I(N__6791));
    Span4Mux_v I__1185 (
            .O(N__6791),
            .I(N__6788));
    Span4Mux_v I__1184 (
            .O(N__6788),
            .I(N__6785));
    Sp12to4 I__1183 (
            .O(N__6785),
            .I(N__6782));
    Span12Mux_h I__1182 (
            .O(N__6782),
            .I(N__6779));
    Odrv12 I__1181 (
            .O(N__6779),
            .I(A_c_6));
    InMux I__1180 (
            .O(N__6776),
            .I(N__6773));
    LocalMux I__1179 (
            .O(N__6773),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ));
    InMux I__1178 (
            .O(N__6770),
            .I(N__6767));
    LocalMux I__1177 (
            .O(N__6767),
            .I(N__6764));
    Span12Mux_v I__1176 (
            .O(N__6764),
            .I(N__6761));
    Span12Mux_h I__1175 (
            .O(N__6761),
            .I(N__6758));
    Span12Mux_v I__1174 (
            .O(N__6758),
            .I(N__6755));
    Odrv12 I__1173 (
            .O(N__6755),
            .I(A_c_2));
    InMux I__1172 (
            .O(N__6752),
            .I(N__6749));
    LocalMux I__1171 (
            .O(N__6749),
            .I(N__6746));
    Odrv4 I__1170 (
            .O(N__6746),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ));
    InMux I__1169 (
            .O(N__6743),
            .I(N__6740));
    LocalMux I__1168 (
            .O(N__6740),
            .I(\U712_REG_SM.STATE_COUNTsr_0 ));
    InMux I__1167 (
            .O(N__6737),
            .I(N__6734));
    LocalMux I__1166 (
            .O(N__6734),
            .I(N__6731));
    Span4Mux_h I__1165 (
            .O(N__6731),
            .I(N__6725));
    InMux I__1164 (
            .O(N__6730),
            .I(N__6722));
    InMux I__1163 (
            .O(N__6729),
            .I(N__6719));
    InMux I__1162 (
            .O(N__6728),
            .I(N__6716));
    Odrv4 I__1161 (
            .O(N__6725),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1160 (
            .O(N__6722),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1159 (
            .O(N__6719),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    LocalMux I__1158 (
            .O(N__6716),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_0 ));
    InMux I__1157 (
            .O(N__6707),
            .I(N__6704));
    LocalMux I__1156 (
            .O(N__6704),
            .I(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ));
    InMux I__1155 (
            .O(N__6701),
            .I(N__6698));
    LocalMux I__1154 (
            .O(N__6698),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_7 ));
    InMux I__1153 (
            .O(N__6695),
            .I(N__6690));
    InMux I__1152 (
            .O(N__6694),
            .I(N__6685));
    InMux I__1151 (
            .O(N__6693),
            .I(N__6685));
    LocalMux I__1150 (
            .O(N__6690),
            .I(\U712_REG_SM.N_307 ));
    LocalMux I__1149 (
            .O(N__6685),
            .I(\U712_REG_SM.N_307 ));
    InMux I__1148 (
            .O(N__6680),
            .I(N__6676));
    InMux I__1147 (
            .O(N__6679),
            .I(N__6673));
    LocalMux I__1146 (
            .O(N__6676),
            .I(\U712_REG_SM.N_553 ));
    LocalMux I__1145 (
            .O(N__6673),
            .I(\U712_REG_SM.N_553 ));
    InMux I__1144 (
            .O(N__6668),
            .I(N__6665));
    LocalMux I__1143 (
            .O(N__6665),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_4 ));
    InMux I__1142 (
            .O(N__6662),
            .I(N__6656));
    InMux I__1141 (
            .O(N__6661),
            .I(N__6656));
    LocalMux I__1140 (
            .O(N__6656),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_5 ));
    InMux I__1139 (
            .O(N__6653),
            .I(N__6650));
    LocalMux I__1138 (
            .O(N__6650),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_6 ));
    IoInMux I__1137 (
            .O(N__6647),
            .I(N__6644));
    LocalMux I__1136 (
            .O(N__6644),
            .I(N__6641));
    IoSpan4Mux I__1135 (
            .O(N__6641),
            .I(N__6638));
    Span4Mux_s3_v I__1134 (
            .O(N__6638),
            .I(N__6635));
    Span4Mux_v I__1133 (
            .O(N__6635),
            .I(N__6632));
    Odrv4 I__1132 (
            .O(N__6632),
            .I(N_130_i));
    InMux I__1131 (
            .O(N__6629),
            .I(N__6626));
    LocalMux I__1130 (
            .O(N__6626),
            .I(N__6623));
    Odrv4 I__1129 (
            .O(N__6623),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ));
    InMux I__1128 (
            .O(N__6620),
            .I(N__6615));
    InMux I__1127 (
            .O(N__6619),
            .I(N__6612));
    InMux I__1126 (
            .O(N__6618),
            .I(N__6609));
    LocalMux I__1125 (
            .O(N__6615),
            .I(N__6606));
    LocalMux I__1124 (
            .O(N__6612),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    LocalMux I__1123 (
            .O(N__6609),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    Odrv4 I__1122 (
            .O(N__6606),
            .I(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ));
    CascadeMux I__1121 (
            .O(N__6599),
            .I(\U712_REG_SM.N_306_cascade_ ));
    CascadeMux I__1120 (
            .O(N__6596),
            .I(\U712_REG_SM.N_399_cascade_ ));
    InMux I__1119 (
            .O(N__6593),
            .I(N__6590));
    LocalMux I__1118 (
            .O(N__6590),
            .I(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ));
    InMux I__1117 (
            .O(N__6587),
            .I(N__6581));
    InMux I__1116 (
            .O(N__6586),
            .I(N__6581));
    LocalMux I__1115 (
            .O(N__6581),
            .I(\U712_REG_SM.N_311 ));
    CascadeMux I__1114 (
            .O(N__6578),
            .I(\U712_REG_SM.N_353_cascade_ ));
    InMux I__1113 (
            .O(N__6575),
            .I(N__6570));
    InMux I__1112 (
            .O(N__6574),
            .I(N__6565));
    InMux I__1111 (
            .O(N__6573),
            .I(N__6565));
    LocalMux I__1110 (
            .O(N__6570),
            .I(N__6562));
    LocalMux I__1109 (
            .O(N__6565),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    Odrv4 I__1108 (
            .O(N__6562),
            .I(\U712_REG_SM.STATE_COUNTZ0Z_2 ));
    InMux I__1107 (
            .O(N__6557),
            .I(N__6554));
    LocalMux I__1106 (
            .O(N__6554),
            .I(N__6551));
    Odrv4 I__1105 (
            .O(N__6551),
            .I(\U712_REG_SM.C3_SYNCZ0Z_0 ));
    InMux I__1104 (
            .O(N__6548),
            .I(N__6545));
    LocalMux I__1103 (
            .O(N__6545),
            .I(\U712_REG_SM.N_322 ));
    InMux I__1102 (
            .O(N__6542),
            .I(N__6535));
    InMux I__1101 (
            .O(N__6541),
            .I(N__6535));
    CascadeMux I__1100 (
            .O(N__6540),
            .I(N__6532));
    LocalMux I__1099 (
            .O(N__6535),
            .I(N__6528));
    InMux I__1098 (
            .O(N__6532),
            .I(N__6525));
    InMux I__1097 (
            .O(N__6531),
            .I(N__6522));
    Span4Mux_h I__1096 (
            .O(N__6528),
            .I(N__6519));
    LocalMux I__1095 (
            .O(N__6525),
            .I(REG_TACK));
    LocalMux I__1094 (
            .O(N__6522),
            .I(REG_TACK));
    Odrv4 I__1093 (
            .O(N__6519),
            .I(REG_TACK));
    CascadeMux I__1092 (
            .O(N__6512),
            .I(\U712_CHIP_RAM.N_356_cascade_ ));
    InMux I__1091 (
            .O(N__6509),
            .I(N__6506));
    LocalMux I__1090 (
            .O(N__6506),
            .I(\U712_CHIP_RAM.N_448 ));
    CascadeMux I__1089 (
            .O(N__6503),
            .I(\U712_CHIP_RAM.N_288_cascade_ ));
    InMux I__1088 (
            .O(N__6500),
            .I(N__6496));
    InMux I__1087 (
            .O(N__6499),
            .I(N__6493));
    LocalMux I__1086 (
            .O(N__6496),
            .I(\U712_CHIP_RAM.N_473 ));
    LocalMux I__1085 (
            .O(N__6493),
            .I(\U712_CHIP_RAM.N_473 ));
    CascadeMux I__1084 (
            .O(N__6488),
            .I(\U712_CHIP_RAM.N_473_cascade_ ));
    InMux I__1083 (
            .O(N__6485),
            .I(N__6482));
    LocalMux I__1082 (
            .O(N__6482),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0 ));
    InMux I__1081 (
            .O(N__6479),
            .I(N__6476));
    LocalMux I__1080 (
            .O(N__6476),
            .I(N__6471));
    InMux I__1079 (
            .O(N__6475),
            .I(N__6466));
    InMux I__1078 (
            .O(N__6474),
            .I(N__6466));
    Odrv4 I__1077 (
            .O(N__6471),
            .I(\U712_CHIP_RAM.N_362 ));
    LocalMux I__1076 (
            .O(N__6466),
            .I(\U712_CHIP_RAM.N_362 ));
    InMux I__1075 (
            .O(N__6461),
            .I(N__6458));
    LocalMux I__1074 (
            .O(N__6458),
            .I(N__6451));
    InMux I__1073 (
            .O(N__6457),
            .I(N__6446));
    InMux I__1072 (
            .O(N__6456),
            .I(N__6446));
    InMux I__1071 (
            .O(N__6455),
            .I(N__6443));
    InMux I__1070 (
            .O(N__6454),
            .I(N__6440));
    Odrv4 I__1069 (
            .O(N__6451),
            .I(\U712_CHIP_RAM.N_463 ));
    LocalMux I__1068 (
            .O(N__6446),
            .I(\U712_CHIP_RAM.N_463 ));
    LocalMux I__1067 (
            .O(N__6443),
            .I(\U712_CHIP_RAM.N_463 ));
    LocalMux I__1066 (
            .O(N__6440),
            .I(\U712_CHIP_RAM.N_463 ));
    CEMux I__1065 (
            .O(N__6431),
            .I(N__6428));
    LocalMux I__1064 (
            .O(N__6428),
            .I(N__6425));
    Odrv4 I__1063 (
            .O(N__6425),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ));
    InMux I__1062 (
            .O(N__6422),
            .I(N__6418));
    InMux I__1061 (
            .O(N__6421),
            .I(N__6415));
    LocalMux I__1060 (
            .O(N__6418),
            .I(N__6410));
    LocalMux I__1059 (
            .O(N__6415),
            .I(N__6410));
    Odrv4 I__1058 (
            .O(N__6410),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ));
    IoInMux I__1057 (
            .O(N__6407),
            .I(N__6404));
    LocalMux I__1056 (
            .O(N__6404),
            .I(N__6401));
    IoSpan4Mux I__1055 (
            .O(N__6401),
            .I(N__6398));
    Span4Mux_s2_v I__1054 (
            .O(N__6398),
            .I(N__6395));
    Sp12to4 I__1053 (
            .O(N__6395),
            .I(N__6392));
    Span12Mux_v I__1052 (
            .O(N__6392),
            .I(N__6388));
    InMux I__1051 (
            .O(N__6391),
            .I(N__6385));
    Odrv12 I__1050 (
            .O(N__6388),
            .I(DBDIR_c));
    LocalMux I__1049 (
            .O(N__6385),
            .I(DBDIR_c));
    CascadeMux I__1048 (
            .O(N__6380),
            .I(N__6377));
    InMux I__1047 (
            .O(N__6377),
            .I(N__6374));
    LocalMux I__1046 (
            .O(N__6374),
            .I(N__6371));
    Odrv4 I__1045 (
            .O(N__6371),
            .I(\U712_CHIP_RAM.N_556 ));
    InMux I__1044 (
            .O(N__6368),
            .I(N__6365));
    LocalMux I__1043 (
            .O(N__6365),
            .I(N__6360));
    InMux I__1042 (
            .O(N__6364),
            .I(N__6357));
    InMux I__1041 (
            .O(N__6363),
            .I(N__6354));
    Odrv4 I__1040 (
            .O(N__6360),
            .I(\U712_CHIP_RAM.N_302 ));
    LocalMux I__1039 (
            .O(N__6357),
            .I(\U712_CHIP_RAM.N_302 ));
    LocalMux I__1038 (
            .O(N__6354),
            .I(\U712_CHIP_RAM.N_302 ));
    InMux I__1037 (
            .O(N__6347),
            .I(N__6344));
    LocalMux I__1036 (
            .O(N__6344),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER19 ));
    CascadeMux I__1035 (
            .O(N__6341),
            .I(\U712_CHIP_RAM.N_355_cascade_ ));
    CascadeMux I__1034 (
            .O(N__6338),
            .I(N__6335));
    InMux I__1033 (
            .O(N__6335),
            .I(N__6332));
    LocalMux I__1032 (
            .O(N__6332),
            .I(N__6329));
    Odrv4 I__1031 (
            .O(N__6329),
            .I(\U712_CHIP_RAM.N_389 ));
    InMux I__1030 (
            .O(N__6326),
            .I(N__6320));
    InMux I__1029 (
            .O(N__6325),
            .I(N__6320));
    LocalMux I__1028 (
            .O(N__6320),
            .I(\U712_CHIP_RAM.N_301 ));
    CascadeMux I__1027 (
            .O(N__6317),
            .I(N__6313));
    CascadeMux I__1026 (
            .O(N__6316),
            .I(N__6309));
    InMux I__1025 (
            .O(N__6313),
            .I(N__6305));
    CascadeMux I__1024 (
            .O(N__6312),
            .I(N__6302));
    InMux I__1023 (
            .O(N__6309),
            .I(N__6298));
    InMux I__1022 (
            .O(N__6308),
            .I(N__6295));
    LocalMux I__1021 (
            .O(N__6305),
            .I(N__6292));
    InMux I__1020 (
            .O(N__6302),
            .I(N__6287));
    InMux I__1019 (
            .O(N__6301),
            .I(N__6287));
    LocalMux I__1018 (
            .O(N__6298),
            .I(\U712_CHIP_RAM.N_289 ));
    LocalMux I__1017 (
            .O(N__6295),
            .I(\U712_CHIP_RAM.N_289 ));
    Odrv4 I__1016 (
            .O(N__6292),
            .I(\U712_CHIP_RAM.N_289 ));
    LocalMux I__1015 (
            .O(N__6287),
            .I(\U712_CHIP_RAM.N_289 ));
    InMux I__1014 (
            .O(N__6278),
            .I(N__6275));
    LocalMux I__1013 (
            .O(N__6275),
            .I(N__6272));
    Odrv4 I__1012 (
            .O(N__6272),
            .I(\U712_CHIP_RAM.N_356 ));
    CascadeMux I__1011 (
            .O(N__6269),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ));
    InMux I__1010 (
            .O(N__6266),
            .I(N__6263));
    LocalMux I__1009 (
            .O(N__6263),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ));
    InMux I__1008 (
            .O(N__6260),
            .I(N__6257));
    LocalMux I__1007 (
            .O(N__6257),
            .I(N__6254));
    Span4Mux_h I__1006 (
            .O(N__6254),
            .I(N__6250));
    InMux I__1005 (
            .O(N__6253),
            .I(N__6247));
    Odrv4 I__1004 (
            .O(N__6250),
            .I(\U712_CHIP_RAM.N_551 ));
    LocalMux I__1003 (
            .O(N__6247),
            .I(\U712_CHIP_RAM.N_551 ));
    CEMux I__1002 (
            .O(N__6242),
            .I(N__6239));
    LocalMux I__1001 (
            .O(N__6239),
            .I(N__6236));
    Span4Mux_v I__1000 (
            .O(N__6236),
            .I(N__6233));
    Odrv4 I__999 (
            .O(N__6233),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0 ));
    InMux I__998 (
            .O(N__6230),
            .I(N__6226));
    InMux I__997 (
            .O(N__6229),
            .I(N__6223));
    LocalMux I__996 (
            .O(N__6226),
            .I(N__6218));
    LocalMux I__995 (
            .O(N__6223),
            .I(N__6218));
    Odrv4 I__994 (
            .O(N__6218),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ));
    InMux I__993 (
            .O(N__6215),
            .I(N__6212));
    LocalMux I__992 (
            .O(N__6212),
            .I(N__6209));
    Span4Mux_v I__991 (
            .O(N__6209),
            .I(N__6206));
    Sp12to4 I__990 (
            .O(N__6206),
            .I(N__6203));
    Span12Mux_h I__989 (
            .O(N__6203),
            .I(N__6200));
    Span12Mux_v I__988 (
            .O(N__6200),
            .I(N__6197));
    Odrv12 I__987 (
            .O(N__6197),
            .I(A_c_20));
    InMux I__986 (
            .O(N__6194),
            .I(N__6190));
    InMux I__985 (
            .O(N__6193),
            .I(N__6187));
    LocalMux I__984 (
            .O(N__6190),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    LocalMux I__983 (
            .O(N__6187),
            .I(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ));
    CascadeMux I__982 (
            .O(N__6182),
            .I(\U712_CHIP_RAM.N_555_cascade_ ));
    InMux I__981 (
            .O(N__6179),
            .I(N__6176));
    LocalMux I__980 (
            .O(N__6176),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16 ));
    InMux I__979 (
            .O(N__6173),
            .I(N__6170));
    LocalMux I__978 (
            .O(N__6170),
            .I(N__6167));
    Odrv4 I__977 (
            .O(N__6167),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0 ));
    CascadeMux I__976 (
            .O(N__6164),
            .I(\U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ));
    CascadeMux I__975 (
            .O(N__6161),
            .I(\U712_REG_SM.N_307_cascade_ ));
    InMux I__974 (
            .O(N__6158),
            .I(N__6153));
    InMux I__973 (
            .O(N__6157),
            .I(N__6150));
    InMux I__972 (
            .O(N__6156),
            .I(N__6147));
    LocalMux I__971 (
            .O(N__6153),
            .I(N__6142));
    LocalMux I__970 (
            .O(N__6150),
            .I(N__6142));
    LocalMux I__969 (
            .O(N__6147),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_3 ));
    Odrv4 I__968 (
            .O(N__6142),
            .I(\U712_REG_SM.STATE_COUNTZ1Z_3 ));
    IoInMux I__967 (
            .O(N__6137),
            .I(N__6134));
    LocalMux I__966 (
            .O(N__6134),
            .I(N__6131));
    Span4Mux_s2_v I__965 (
            .O(N__6131),
            .I(N__6128));
    Sp12to4 I__964 (
            .O(N__6128),
            .I(N__6125));
    Span12Mux_h I__963 (
            .O(N__6125),
            .I(N__6120));
    InMux I__962 (
            .O(N__6124),
            .I(N__6117));
    InMux I__961 (
            .O(N__6123),
            .I(N__6114));
    Odrv12 I__960 (
            .O(N__6120),
            .I(REGENn_c));
    LocalMux I__959 (
            .O(N__6117),
            .I(REGENn_c));
    LocalMux I__958 (
            .O(N__6114),
            .I(REGENn_c));
    InMux I__957 (
            .O(N__6107),
            .I(N__6104));
    LocalMux I__956 (
            .O(N__6104),
            .I(\U712_REG_SM.REGENn_e_1 ));
    InMux I__955 (
            .O(N__6101),
            .I(N__6095));
    InMux I__954 (
            .O(N__6100),
            .I(N__6095));
    LocalMux I__953 (
            .O(N__6095),
            .I(N__6090));
    InMux I__952 (
            .O(N__6094),
            .I(N__6087));
    InMux I__951 (
            .O(N__6093),
            .I(N__6084));
    Odrv4 I__950 (
            .O(N__6090),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__949 (
            .O(N__6087),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    LocalMux I__948 (
            .O(N__6084),
            .I(\U712_REG_SM.REG_CYCLE_STARTZ0 ));
    InMux I__947 (
            .O(N__6077),
            .I(N__6070));
    InMux I__946 (
            .O(N__6076),
            .I(N__6070));
    InMux I__945 (
            .O(N__6075),
            .I(N__6067));
    LocalMux I__944 (
            .O(N__6070),
            .I(N__6064));
    LocalMux I__943 (
            .O(N__6067),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    Odrv4 I__942 (
            .O(N__6064),
            .I(\U712_REG_SM.WRITE_CYCLEZ0 ));
    InMux I__941 (
            .O(N__6059),
            .I(N__6056));
    LocalMux I__940 (
            .O(N__6056),
            .I(N__6053));
    Span12Mux_h I__939 (
            .O(N__6053),
            .I(N__6050));
    Odrv12 I__938 (
            .O(N__6050),
            .I(A_c_12));
    IoInMux I__937 (
            .O(N__6047),
            .I(N__6044));
    LocalMux I__936 (
            .O(N__6044),
            .I(N__6041));
    IoSpan4Mux I__935 (
            .O(N__6041),
            .I(N__6038));
    Span4Mux_s2_v I__934 (
            .O(N__6038),
            .I(N__6034));
    InMux I__933 (
            .O(N__6037),
            .I(N__6031));
    Sp12to4 I__932 (
            .O(N__6034),
            .I(N__6028));
    LocalMux I__931 (
            .O(N__6031),
            .I(N__6025));
    Span12Mux_s8_v I__930 (
            .O(N__6028),
            .I(N__6022));
    Span4Mux_v I__929 (
            .O(N__6025),
            .I(N__6019));
    Span12Mux_v I__928 (
            .O(N__6022),
            .I(N__6016));
    Sp12to4 I__927 (
            .O(N__6019),
            .I(N__6013));
    Span12Mux_h I__926 (
            .O(N__6016),
            .I(N__6010));
    Span12Mux_h I__925 (
            .O(N__6013),
            .I(N__6007));
    Odrv12 I__924 (
            .O(N__6010),
            .I(A_c_11));
    Odrv12 I__923 (
            .O(N__6007),
            .I(A_c_11));
    InMux I__922 (
            .O(N__6002),
            .I(N__5998));
    InMux I__921 (
            .O(N__6001),
            .I(N__5995));
    LocalMux I__920 (
            .O(N__5998),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    LocalMux I__919 (
            .O(N__5995),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ));
    CascadeMux I__918 (
            .O(N__5990),
            .I(N__5987));
    InMux I__917 (
            .O(N__5987),
            .I(N__5984));
    LocalMux I__916 (
            .O(N__5984),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ));
    InMux I__915 (
            .O(N__5981),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ));
    InMux I__914 (
            .O(N__5978),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ));
    CascadeMux I__913 (
            .O(N__5975),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ));
    InMux I__912 (
            .O(N__5972),
            .I(N__5968));
    InMux I__911 (
            .O(N__5971),
            .I(N__5965));
    LocalMux I__910 (
            .O(N__5968),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    LocalMux I__909 (
            .O(N__5965),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ));
    InMux I__908 (
            .O(N__5960),
            .I(N__5957));
    LocalMux I__907 (
            .O(N__5957),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ));
    InMux I__906 (
            .O(N__5954),
            .I(N__5950));
    InMux I__905 (
            .O(N__5953),
            .I(N__5947));
    LocalMux I__904 (
            .O(N__5950),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ));
    LocalMux I__903 (
            .O(N__5947),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ));
    InMux I__902 (
            .O(N__5942),
            .I(N__5931));
    InMux I__901 (
            .O(N__5941),
            .I(N__5931));
    InMux I__900 (
            .O(N__5940),
            .I(N__5924));
    InMux I__899 (
            .O(N__5939),
            .I(N__5924));
    InMux I__898 (
            .O(N__5938),
            .I(N__5924));
    InMux I__897 (
            .O(N__5937),
            .I(N__5919));
    InMux I__896 (
            .O(N__5936),
            .I(N__5919));
    LocalMux I__895 (
            .O(N__5931),
            .I(N__5916));
    LocalMux I__894 (
            .O(N__5924),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    LocalMux I__893 (
            .O(N__5919),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    Odrv4 I__892 (
            .O(N__5916),
            .I(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ));
    CascadeMux I__891 (
            .O(N__5909),
            .I(N__5906));
    InMux I__890 (
            .O(N__5906),
            .I(N__5903));
    LocalMux I__889 (
            .O(N__5903),
            .I(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ));
    CascadeMux I__888 (
            .O(N__5900),
            .I(N__5897));
    InMux I__887 (
            .O(N__5897),
            .I(N__5893));
    InMux I__886 (
            .O(N__5896),
            .I(N__5890));
    LocalMux I__885 (
            .O(N__5893),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    LocalMux I__884 (
            .O(N__5890),
            .I(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ));
    CascadeMux I__883 (
            .O(N__5885),
            .I(N__5882));
    InMux I__882 (
            .O(N__5882),
            .I(N__5875));
    InMux I__881 (
            .O(N__5881),
            .I(N__5875));
    InMux I__880 (
            .O(N__5880),
            .I(N__5872));
    LocalMux I__879 (
            .O(N__5875),
            .I(N__5866));
    LocalMux I__878 (
            .O(N__5872),
            .I(N__5866));
    InMux I__877 (
            .O(N__5871),
            .I(N__5863));
    Span4Mux_v I__876 (
            .O(N__5866),
            .I(N__5860));
    LocalMux I__875 (
            .O(N__5863),
            .I(CPU_TACKm));
    Odrv4 I__874 (
            .O(N__5860),
            .I(CPU_TACKm));
    InMux I__873 (
            .O(N__5855),
            .I(N__5852));
    LocalMux I__872 (
            .O(N__5852),
            .I(\U712_CYCLE_TERM.TACK_EN6_0 ));
    CascadeMux I__871 (
            .O(N__5849),
            .I(N__5842));
    CascadeMux I__870 (
            .O(N__5848),
            .I(N__5838));
    InMux I__869 (
            .O(N__5847),
            .I(N__5834));
    InMux I__868 (
            .O(N__5846),
            .I(N__5827));
    InMux I__867 (
            .O(N__5845),
            .I(N__5827));
    InMux I__866 (
            .O(N__5842),
            .I(N__5827));
    InMux I__865 (
            .O(N__5841),
            .I(N__5820));
    InMux I__864 (
            .O(N__5838),
            .I(N__5820));
    InMux I__863 (
            .O(N__5837),
            .I(N__5820));
    LocalMux I__862 (
            .O(N__5834),
            .I(N__5815));
    LocalMux I__861 (
            .O(N__5827),
            .I(N__5810));
    LocalMux I__860 (
            .O(N__5820),
            .I(N__5810));
    InMux I__859 (
            .O(N__5819),
            .I(N__5805));
    InMux I__858 (
            .O(N__5818),
            .I(N__5805));
    Odrv12 I__857 (
            .O(N__5815),
            .I(DBR_SYNCZ0Z_1));
    Odrv4 I__856 (
            .O(N__5810),
            .I(DBR_SYNCZ0Z_1));
    LocalMux I__855 (
            .O(N__5805),
            .I(DBR_SYNCZ0Z_1));
    CascadeMux I__854 (
            .O(N__5798),
            .I(N__5794));
    InMux I__853 (
            .O(N__5797),
            .I(N__5791));
    InMux I__852 (
            .O(N__5794),
            .I(N__5788));
    LocalMux I__851 (
            .O(N__5791),
            .I(DBR_SYNC_i_1));
    LocalMux I__850 (
            .O(N__5788),
            .I(DBR_SYNC_i_1));
    InMux I__849 (
            .O(N__5783),
            .I(N__5780));
    LocalMux I__848 (
            .O(N__5780),
            .I(\U712_CHIP_RAM.N_360 ));
    InMux I__847 (
            .O(N__5777),
            .I(N__5773));
    InMux I__846 (
            .O(N__5776),
            .I(N__5770));
    LocalMux I__845 (
            .O(N__5773),
            .I(\U712_CHIP_RAM.N_418 ));
    LocalMux I__844 (
            .O(N__5770),
            .I(\U712_CHIP_RAM.N_418 ));
    InMux I__843 (
            .O(N__5765),
            .I(N__5762));
    LocalMux I__842 (
            .O(N__5762),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0 ));
    CascadeMux I__841 (
            .O(N__5759),
            .I(\U712_REG_SM.N_400_cascade_ ));
    CascadeMux I__840 (
            .O(N__5756),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ));
    CascadeMux I__839 (
            .O(N__5753),
            .I(N__5750));
    InMux I__838 (
            .O(N__5750),
            .I(N__5747));
    LocalMux I__837 (
            .O(N__5747),
            .I(\U712_CHIP_RAM.N_405 ));
    InMux I__836 (
            .O(N__5744),
            .I(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ));
    CascadeMux I__835 (
            .O(N__5741),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ));
    InMux I__834 (
            .O(N__5738),
            .I(N__5735));
    LocalMux I__833 (
            .O(N__5735),
            .I(N__5732));
    Odrv4 I__832 (
            .O(N__5732),
            .I(\U712_CHIP_RAM.N_439 ));
    InMux I__831 (
            .O(N__5729),
            .I(N__5726));
    LocalMux I__830 (
            .O(N__5726),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0 ));
    CascadeMux I__829 (
            .O(N__5723),
            .I(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ));
    CascadeMux I__828 (
            .O(N__5720),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ));
    IoInMux I__827 (
            .O(N__5717),
            .I(N__5714));
    LocalMux I__826 (
            .O(N__5714),
            .I(N__5711));
    Span4Mux_s2_h I__825 (
            .O(N__5711),
            .I(N__5708));
    Span4Mux_h I__824 (
            .O(N__5708),
            .I(N__5705));
    Sp12to4 I__823 (
            .O(N__5705),
            .I(N__5702));
    Span12Mux_s11_v I__822 (
            .O(N__5702),
            .I(N__5699));
    Span12Mux_h I__821 (
            .O(N__5699),
            .I(N__5696));
    Odrv12 I__820 (
            .O(N__5696),
            .I(CLK_EN_c));
    CEMux I__819 (
            .O(N__5693),
            .I(N__5690));
    LocalMux I__818 (
            .O(N__5690),
            .I(N__5687));
    Span4Mux_h I__817 (
            .O(N__5687),
            .I(N__5684));
    Odrv4 I__816 (
            .O(N__5684),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ));
    CascadeMux I__815 (
            .O(N__5681),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_ ));
    InMux I__814 (
            .O(N__5678),
            .I(N__5675));
    LocalMux I__813 (
            .O(N__5675),
            .I(N__5672));
    Span4Mux_v I__812 (
            .O(N__5672),
            .I(N__5664));
    InMux I__811 (
            .O(N__5671),
            .I(N__5661));
    InMux I__810 (
            .O(N__5670),
            .I(N__5656));
    InMux I__809 (
            .O(N__5669),
            .I(N__5656));
    InMux I__808 (
            .O(N__5668),
            .I(N__5653));
    InMux I__807 (
            .O(N__5667),
            .I(N__5650));
    Odrv4 I__806 (
            .O(N__5664),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__805 (
            .O(N__5661),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__804 (
            .O(N__5656),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__803 (
            .O(N__5653),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    LocalMux I__802 (
            .O(N__5650),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ));
    InMux I__801 (
            .O(N__5639),
            .I(N__5633));
    InMux I__800 (
            .O(N__5638),
            .I(N__5626));
    InMux I__799 (
            .O(N__5637),
            .I(N__5626));
    InMux I__798 (
            .O(N__5636),
            .I(N__5626));
    LocalMux I__797 (
            .O(N__5633),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ));
    LocalMux I__796 (
            .O(N__5626),
            .I(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ));
    CascadeMux I__795 (
            .O(N__5621),
            .I(N__5618));
    InMux I__794 (
            .O(N__5618),
            .I(N__5615));
    LocalMux I__793 (
            .O(N__5615),
            .I(\U712_CHIP_RAM.N_445 ));
    CascadeMux I__792 (
            .O(N__5612),
            .I(N__5609));
    InMux I__791 (
            .O(N__5609),
            .I(N__5606));
    LocalMux I__790 (
            .O(N__5606),
            .I(\U712_CHIP_RAM.N_208 ));
    InMux I__789 (
            .O(N__5603),
            .I(N__5599));
    InMux I__788 (
            .O(N__5602),
            .I(N__5596));
    LocalMux I__787 (
            .O(N__5599),
            .I(\U712_CHIP_RAM.N_303 ));
    LocalMux I__786 (
            .O(N__5596),
            .I(\U712_CHIP_RAM.N_303 ));
    CascadeMux I__785 (
            .O(N__5591),
            .I(\U712_CHIP_RAM.N_443_cascade_ ));
    InMux I__784 (
            .O(N__5588),
            .I(N__5585));
    LocalMux I__783 (
            .O(N__5585),
            .I(\U712_CHIP_RAM.N_204 ));
    CascadeMux I__782 (
            .O(N__5582),
            .I(\U712_CHIP_RAM.N_463_cascade_ ));
    CascadeMux I__781 (
            .O(N__5579),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ));
    CascadeMux I__780 (
            .O(N__5576),
            .I(N__5573));
    InMux I__779 (
            .O(N__5573),
            .I(N__5570));
    LocalMux I__778 (
            .O(N__5570),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ));
    InMux I__777 (
            .O(N__5567),
            .I(N__5564));
    LocalMux I__776 (
            .O(N__5564),
            .I(N__5561));
    Span4Mux_v I__775 (
            .O(N__5561),
            .I(N__5558));
    Span4Mux_v I__774 (
            .O(N__5558),
            .I(N__5555));
    Sp12to4 I__773 (
            .O(N__5555),
            .I(N__5552));
    Span12Mux_h I__772 (
            .O(N__5552),
            .I(N__5549));
    Odrv12 I__771 (
            .O(N__5549),
            .I(A_c_17));
    CascadeMux I__770 (
            .O(N__5546),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ));
    InMux I__769 (
            .O(N__5543),
            .I(N__5540));
    LocalMux I__768 (
            .O(N__5540),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ));
    InMux I__767 (
            .O(N__5537),
            .I(N__5534));
    LocalMux I__766 (
            .O(N__5534),
            .I(N__5531));
    Span4Mux_v I__765 (
            .O(N__5531),
            .I(N__5528));
    Odrv4 I__764 (
            .O(N__5528),
            .I(\U712_CHIP_RAM.N_346 ));
    InMux I__763 (
            .O(N__5525),
            .I(N__5520));
    InMux I__762 (
            .O(N__5524),
            .I(N__5515));
    InMux I__761 (
            .O(N__5523),
            .I(N__5515));
    LocalMux I__760 (
            .O(N__5520),
            .I(\U712_CHIP_RAM.N_388 ));
    LocalMux I__759 (
            .O(N__5515),
            .I(\U712_CHIP_RAM.N_388 ));
    InMux I__758 (
            .O(N__5510),
            .I(N__5505));
    CascadeMux I__757 (
            .O(N__5509),
            .I(N__5501));
    InMux I__756 (
            .O(N__5508),
            .I(N__5498));
    LocalMux I__755 (
            .O(N__5505),
            .I(N__5495));
    CascadeMux I__754 (
            .O(N__5504),
            .I(N__5492));
    InMux I__753 (
            .O(N__5501),
            .I(N__5488));
    LocalMux I__752 (
            .O(N__5498),
            .I(N__5483));
    Span4Mux_v I__751 (
            .O(N__5495),
            .I(N__5483));
    InMux I__750 (
            .O(N__5492),
            .I(N__5480));
    InMux I__749 (
            .O(N__5491),
            .I(N__5477));
    LocalMux I__748 (
            .O(N__5488),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    Odrv4 I__747 (
            .O(N__5483),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__746 (
            .O(N__5480),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    LocalMux I__745 (
            .O(N__5477),
            .I(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ));
    SRMux I__744 (
            .O(N__5468),
            .I(N__5465));
    LocalMux I__743 (
            .O(N__5465),
            .I(N__5461));
    InMux I__742 (
            .O(N__5464),
            .I(N__5458));
    Span4Mux_h I__741 (
            .O(N__5461),
            .I(N__5455));
    LocalMux I__740 (
            .O(N__5458),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    Odrv4 I__739 (
            .O(N__5455),
            .I(\U712_CHIP_RAM.REFRESH_RST ));
    CascadeMux I__738 (
            .O(N__5450),
            .I(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ));
    InMux I__737 (
            .O(N__5447),
            .I(N__5443));
    InMux I__736 (
            .O(N__5446),
            .I(N__5440));
    LocalMux I__735 (
            .O(N__5443),
            .I(\U712_REG_SM.START_RSTZ0 ));
    LocalMux I__734 (
            .O(N__5440),
            .I(\U712_REG_SM.START_RSTZ0 ));
    InMux I__733 (
            .O(N__5435),
            .I(N__5431));
    IoInMux I__732 (
            .O(N__5434),
            .I(N__5428));
    LocalMux I__731 (
            .O(N__5431),
            .I(N__5425));
    LocalMux I__730 (
            .O(N__5428),
            .I(N__5422));
    Span4Mux_v I__729 (
            .O(N__5425),
            .I(N__5419));
    IoSpan4Mux I__728 (
            .O(N__5422),
            .I(N__5416));
    Sp12to4 I__727 (
            .O(N__5419),
            .I(N__5413));
    IoSpan4Mux I__726 (
            .O(N__5416),
            .I(N__5410));
    Span12Mux_h I__725 (
            .O(N__5413),
            .I(N__5407));
    IoSpan4Mux I__724 (
            .O(N__5410),
            .I(N__5404));
    Odrv12 I__723 (
            .O(N__5407),
            .I(C1_c));
    Odrv4 I__722 (
            .O(N__5404),
            .I(C1_c));
    InMux I__721 (
            .O(N__5399),
            .I(N__5396));
    LocalMux I__720 (
            .O(N__5396),
            .I(\U712_REG_SM.C1_SYNCZ0Z_0 ));
    IoInMux I__719 (
            .O(N__5393),
            .I(N__5390));
    LocalMux I__718 (
            .O(N__5390),
            .I(N__5387));
    IoSpan4Mux I__717 (
            .O(N__5387),
            .I(N__5384));
    Span4Mux_s2_v I__716 (
            .O(N__5384),
            .I(N__5381));
    Span4Mux_v I__715 (
            .O(N__5381),
            .I(N__5378));
    Span4Mux_h I__714 (
            .O(N__5378),
            .I(N__5375));
    Odrv4 I__713 (
            .O(N__5375),
            .I(CRCSn_c));
    IoInMux I__712 (
            .O(N__5372),
            .I(N__5369));
    LocalMux I__711 (
            .O(N__5369),
            .I(N__5366));
    IoSpan4Mux I__710 (
            .O(N__5366),
            .I(N__5363));
    Sp12to4 I__709 (
            .O(N__5363),
            .I(N__5360));
    Span12Mux_s9_v I__708 (
            .O(N__5360),
            .I(N__5357));
    Odrv12 I__707 (
            .O(N__5357),
            .I(RASn_c));
    IoInMux I__706 (
            .O(N__5354),
            .I(N__5351));
    LocalMux I__705 (
            .O(N__5351),
            .I(N__5348));
    Span12Mux_s10_v I__704 (
            .O(N__5348),
            .I(N__5345));
    Odrv12 I__703 (
            .O(N__5345),
            .I(CMA_c_0));
    IoInMux I__702 (
            .O(N__5342),
            .I(N__5339));
    LocalMux I__701 (
            .O(N__5339),
            .I(N__5336));
    Span12Mux_s10_v I__700 (
            .O(N__5336),
            .I(N__5333));
    Odrv12 I__699 (
            .O(N__5333),
            .I(CMA_c_10));
    IoInMux I__698 (
            .O(N__5330),
            .I(N__5327));
    LocalMux I__697 (
            .O(N__5327),
            .I(N__5324));
    Span12Mux_s10_v I__696 (
            .O(N__5324),
            .I(N__5321));
    Odrv12 I__695 (
            .O(N__5321),
            .I(CMA_c_2));
    IoInMux I__694 (
            .O(N__5318),
            .I(N__5314));
    InMux I__693 (
            .O(N__5317),
            .I(N__5311));
    LocalMux I__692 (
            .O(N__5314),
            .I(N__5308));
    LocalMux I__691 (
            .O(N__5311),
            .I(N__5305));
    Span12Mux_s4_v I__690 (
            .O(N__5308),
            .I(N__5302));
    Span4Mux_h I__689 (
            .O(N__5305),
            .I(N__5299));
    Span12Mux_v I__688 (
            .O(N__5302),
            .I(N__5296));
    Span4Mux_v I__687 (
            .O(N__5299),
            .I(N__5293));
    Span12Mux_h I__686 (
            .O(N__5296),
            .I(N__5290));
    Sp12to4 I__685 (
            .O(N__5293),
            .I(N__5287));
    Odrv12 I__684 (
            .O(N__5290),
            .I(A_c_9));
    Odrv12 I__683 (
            .O(N__5287),
            .I(A_c_9));
    InMux I__682 (
            .O(N__5282),
            .I(N__5279));
    LocalMux I__681 (
            .O(N__5279),
            .I(\U712_CYCLE_TERM.N_312 ));
    InMux I__680 (
            .O(N__5276),
            .I(N__5270));
    InMux I__679 (
            .O(N__5275),
            .I(N__5270));
    LocalMux I__678 (
            .O(N__5270),
            .I(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ));
    InMux I__677 (
            .O(N__5267),
            .I(N__5262));
    InMux I__676 (
            .O(N__5266),
            .I(N__5257));
    InMux I__675 (
            .O(N__5265),
            .I(N__5257));
    LocalMux I__674 (
            .O(N__5262),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    LocalMux I__673 (
            .O(N__5257),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ));
    IoInMux I__672 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__671 (
            .O(N__5249),
            .I(N__5245));
    IoInMux I__670 (
            .O(N__5248),
            .I(N__5242));
    IoSpan4Mux I__669 (
            .O(N__5245),
            .I(N__5238));
    LocalMux I__668 (
            .O(N__5242),
            .I(N__5235));
    IoInMux I__667 (
            .O(N__5241),
            .I(N__5232));
    Sp12to4 I__666 (
            .O(N__5238),
            .I(N__5229));
    Span4Mux_s3_v I__665 (
            .O(N__5235),
            .I(N__5226));
    LocalMux I__664 (
            .O(N__5232),
            .I(N__5223));
    Span12Mux_s7_h I__663 (
            .O(N__5229),
            .I(N__5220));
    Sp12to4 I__662 (
            .O(N__5226),
            .I(N__5217));
    IoSpan4Mux I__661 (
            .O(N__5223),
            .I(N__5214));
    Span12Mux_h I__660 (
            .O(N__5220),
            .I(N__5209));
    Span12Mux_h I__659 (
            .O(N__5217),
            .I(N__5209));
    Sp12to4 I__658 (
            .O(N__5214),
            .I(N__5206));
    Span12Mux_v I__657 (
            .O(N__5209),
            .I(N__5200));
    Span12Mux_h I__656 (
            .O(N__5206),
            .I(N__5200));
    InMux I__655 (
            .O(N__5205),
            .I(N__5197));
    Odrv12 I__654 (
            .O(N__5200),
            .I(TACK_OUTn));
    LocalMux I__653 (
            .O(N__5197),
            .I(TACK_OUTn));
    InMux I__652 (
            .O(N__5192),
            .I(N__5189));
    LocalMux I__651 (
            .O(N__5189),
            .I(N__5185));
    InMux I__650 (
            .O(N__5188),
            .I(N__5182));
    Span4Mux_v I__649 (
            .O(N__5185),
            .I(N__5179));
    LocalMux I__648 (
            .O(N__5182),
            .I(N__5176));
    Span4Mux_h I__647 (
            .O(N__5179),
            .I(N__5171));
    Span4Mux_v I__646 (
            .O(N__5176),
            .I(N__5171));
    Span4Mux_h I__645 (
            .O(N__5171),
            .I(N__5168));
    Sp12to4 I__644 (
            .O(N__5168),
            .I(N__5165));
    Odrv12 I__643 (
            .O(N__5165),
            .I(DBRn_c));
    InMux I__642 (
            .O(N__5162),
            .I(N__5159));
    LocalMux I__641 (
            .O(N__5159),
            .I(DBR_SYNCZ0Z_0));
    InMux I__640 (
            .O(N__5156),
            .I(N__5152));
    InMux I__639 (
            .O(N__5155),
            .I(N__5149));
    LocalMux I__638 (
            .O(N__5152),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    LocalMux I__637 (
            .O(N__5149),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ));
    InMux I__636 (
            .O(N__5144),
            .I(N__5136));
    InMux I__635 (
            .O(N__5143),
            .I(N__5136));
    InMux I__634 (
            .O(N__5142),
            .I(N__5131));
    InMux I__633 (
            .O(N__5141),
            .I(N__5131));
    LocalMux I__632 (
            .O(N__5136),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    LocalMux I__631 (
            .O(N__5131),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ));
    CascadeMux I__630 (
            .O(N__5126),
            .I(N__5123));
    InMux I__629 (
            .O(N__5123),
            .I(N__5120));
    LocalMux I__628 (
            .O(N__5120),
            .I(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ));
    InMux I__627 (
            .O(N__5117),
            .I(N__5108));
    InMux I__626 (
            .O(N__5116),
            .I(N__5108));
    InMux I__625 (
            .O(N__5115),
            .I(N__5108));
    LocalMux I__624 (
            .O(N__5108),
            .I(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ));
    IoInMux I__623 (
            .O(N__5105),
            .I(N__5102));
    LocalMux I__622 (
            .O(N__5102),
            .I(N__5099));
    IoSpan4Mux I__621 (
            .O(N__5099),
            .I(N__5096));
    Span4Mux_s3_h I__620 (
            .O(N__5096),
            .I(N__5093));
    Span4Mux_v I__619 (
            .O(N__5093),
            .I(N__5089));
    InMux I__618 (
            .O(N__5092),
            .I(N__5086));
    Span4Mux_h I__617 (
            .O(N__5089),
            .I(N__5083));
    LocalMux I__616 (
            .O(N__5086),
            .I(N__5080));
    Sp12to4 I__615 (
            .O(N__5083),
            .I(N__5077));
    Span4Mux_v I__614 (
            .O(N__5080),
            .I(N__5074));
    Span12Mux_h I__613 (
            .O(N__5077),
            .I(N__5069));
    Sp12to4 I__612 (
            .O(N__5074),
            .I(N__5069));
    Span12Mux_h I__611 (
            .O(N__5069),
            .I(N__5066));
    Odrv12 I__610 (
            .O(N__5066),
            .I(C3_c));
    InMux I__609 (
            .O(N__5063),
            .I(N__5060));
    LocalMux I__608 (
            .O(N__5060),
            .I(N__5056));
    InMux I__607 (
            .O(N__5059),
            .I(N__5053));
    Odrv12 I__606 (
            .O(N__5056),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    LocalMux I__605 (
            .O(N__5053),
            .I(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ));
    IoInMux I__604 (
            .O(N__5048),
            .I(N__5045));
    LocalMux I__603 (
            .O(N__5045),
            .I(N__5042));
    Span4Mux_s3_v I__602 (
            .O(N__5042),
            .I(N__5039));
    Span4Mux_h I__601 (
            .O(N__5039),
            .I(N__5036));
    Span4Mux_v I__600 (
            .O(N__5036),
            .I(N__5033));
    Span4Mux_v I__599 (
            .O(N__5033),
            .I(N__5030));
    Span4Mux_v I__598 (
            .O(N__5030),
            .I(N__5026));
    InMux I__597 (
            .O(N__5029),
            .I(N__5023));
    Odrv4 I__596 (
            .O(N__5026),
            .I(LATCH_CLK_c));
    LocalMux I__595 (
            .O(N__5023),
            .I(LATCH_CLK_c));
    InMux I__594 (
            .O(N__5018),
            .I(N__5015));
    LocalMux I__593 (
            .O(N__5015),
            .I(N__5012));
    Span4Mux_h I__592 (
            .O(N__5012),
            .I(N__5008));
    InMux I__591 (
            .O(N__5011),
            .I(N__5005));
    Span4Mux_h I__590 (
            .O(N__5008),
            .I(N__5000));
    LocalMux I__589 (
            .O(N__5005),
            .I(N__5000));
    Span4Mux_v I__588 (
            .O(N__5000),
            .I(N__4997));
    Sp12to4 I__587 (
            .O(N__4997),
            .I(N__4994));
    Span12Mux_h I__586 (
            .O(N__4994),
            .I(N__4991));
    Span12Mux_v I__585 (
            .O(N__4991),
            .I(N__4988));
    Odrv12 I__584 (
            .O(N__4988),
            .I(TSn_c));
    CascadeMux I__583 (
            .O(N__4985),
            .I(N__4982));
    InMux I__582 (
            .O(N__4982),
            .I(N__4979));
    LocalMux I__581 (
            .O(N__4979),
            .I(N__4976));
    Span4Mux_v I__580 (
            .O(N__4976),
            .I(N__4973));
    Sp12to4 I__579 (
            .O(N__4973),
            .I(N__4970));
    Span12Mux_h I__578 (
            .O(N__4970),
            .I(N__4967));
    Span12Mux_v I__577 (
            .O(N__4967),
            .I(N__4964));
    Odrv12 I__576 (
            .O(N__4964),
            .I(REGSPACEn_c));
    InMux I__575 (
            .O(N__4961),
            .I(N__4958));
    LocalMux I__574 (
            .O(N__4958),
            .I(\U712_REG_SM.N_414 ));
    CascadeMux I__573 (
            .O(N__4955),
            .I(\U712_CYCLE_TERM.N_452_cascade_ ));
    InMux I__572 (
            .O(N__4952),
            .I(N__4949));
    LocalMux I__571 (
            .O(N__4949),
            .I(N__4946));
    Span12Mux_h I__570 (
            .O(N__4946),
            .I(N__4943));
    Span12Mux_v I__569 (
            .O(N__4943),
            .I(N__4940));
    Odrv12 I__568 (
            .O(N__4940),
            .I(RAMSPACEn_c));
    CascadeMux I__567 (
            .O(N__4937),
            .I(\U712_CHIP_RAM.N_417_cascade_ ));
    InMux I__566 (
            .O(N__4934),
            .I(N__4929));
    InMux I__565 (
            .O(N__4933),
            .I(N__4924));
    InMux I__564 (
            .O(N__4932),
            .I(N__4924));
    LocalMux I__563 (
            .O(N__4929),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    LocalMux I__562 (
            .O(N__4924),
            .I(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ));
    CascadeMux I__561 (
            .O(N__4919),
            .I(N__4916));
    InMux I__560 (
            .O(N__4916),
            .I(N__4913));
    LocalMux I__559 (
            .O(N__4913),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ));
    InMux I__558 (
            .O(N__4910),
            .I(N__4907));
    LocalMux I__557 (
            .O(N__4907),
            .I(\U712_CHIP_RAM.N_206 ));
    InMux I__556 (
            .O(N__4904),
            .I(N__4901));
    LocalMux I__555 (
            .O(N__4901),
            .I(\U712_CHIP_RAM.N_457 ));
    InMux I__554 (
            .O(N__4898),
            .I(N__4895));
    LocalMux I__553 (
            .O(N__4895),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ));
    InMux I__552 (
            .O(N__4892),
            .I(N__4886));
    InMux I__551 (
            .O(N__4891),
            .I(N__4886));
    LocalMux I__550 (
            .O(N__4886),
            .I(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ));
    InMux I__549 (
            .O(N__4883),
            .I(N__4880));
    LocalMux I__548 (
            .O(N__4880),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1 ));
    InMux I__547 (
            .O(N__4877),
            .I(N__4874));
    LocalMux I__546 (
            .O(N__4874),
            .I(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0 ));
    CascadeMux I__545 (
            .O(N__4871),
            .I(\U712_CHIP_RAM.N_556_cascade_ ));
    InMux I__544 (
            .O(N__4868),
            .I(N__4865));
    LocalMux I__543 (
            .O(N__4865),
            .I(\U712_CHIP_RAM.N_202 ));
    CascadeMux I__542 (
            .O(N__4862),
            .I(\U712_CHIP_RAM.N_388_cascade_ ));
    InMux I__541 (
            .O(N__4859),
            .I(N__4856));
    LocalMux I__540 (
            .O(N__4856),
            .I(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0 ));
    InMux I__539 (
            .O(N__4853),
            .I(N__4849));
    InMux I__538 (
            .O(N__4852),
            .I(N__4846));
    LocalMux I__537 (
            .O(N__4849),
            .I(N__4843));
    LocalMux I__536 (
            .O(N__4846),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    Odrv12 I__535 (
            .O(N__4843),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ));
    InMux I__534 (
            .O(N__4838),
            .I(N__4835));
    LocalMux I__533 (
            .O(N__4835),
            .I(N__4832));
    Odrv4 I__532 (
            .O(N__4832),
            .I(\U712_CHIP_RAM.REFRESH5lto7_0 ));
    InMux I__531 (
            .O(N__4829),
            .I(N__4826));
    LocalMux I__530 (
            .O(N__4826),
            .I(N__4823));
    Odrv12 I__529 (
            .O(N__4823),
            .I(\U712_CHIP_RAM.REFRESH5lt7 ));
    CascadeMux I__528 (
            .O(N__4820),
            .I(N__4816));
    InMux I__527 (
            .O(N__4819),
            .I(N__4810));
    InMux I__526 (
            .O(N__4816),
            .I(N__4810));
    InMux I__525 (
            .O(N__4815),
            .I(N__4807));
    LocalMux I__524 (
            .O(N__4810),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    LocalMux I__523 (
            .O(N__4807),
            .I(\U712_CHIP_RAM.REFRESHZ0 ));
    CascadeMux I__522 (
            .O(N__4802),
            .I(N__4798));
    InMux I__521 (
            .O(N__4801),
            .I(N__4795));
    InMux I__520 (
            .O(N__4798),
            .I(N__4792));
    LocalMux I__519 (
            .O(N__4795),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    LocalMux I__518 (
            .O(N__4792),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ));
    InMux I__517 (
            .O(N__4787),
            .I(N__4783));
    InMux I__516 (
            .O(N__4786),
            .I(N__4780));
    LocalMux I__515 (
            .O(N__4783),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    LocalMux I__514 (
            .O(N__4780),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ));
    InMux I__513 (
            .O(N__4775),
            .I(N__4772));
    LocalMux I__512 (
            .O(N__4772),
            .I(N__4769));
    Sp12to4 I__511 (
            .O(N__4769),
            .I(N__4766));
    Span12Mux_v I__510 (
            .O(N__4766),
            .I(N__4763));
    Span12Mux_h I__509 (
            .O(N__4763),
            .I(N__4760));
    Odrv12 I__508 (
            .O(N__4760),
            .I(A_c_16));
    CascadeMux I__507 (
            .O(N__4757),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ));
    InMux I__506 (
            .O(N__4754),
            .I(N__4750));
    InMux I__505 (
            .O(N__4753),
            .I(N__4747));
    LocalMux I__504 (
            .O(N__4750),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    LocalMux I__503 (
            .O(N__4747),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ));
    InMux I__502 (
            .O(N__4742),
            .I(N__4738));
    InMux I__501 (
            .O(N__4741),
            .I(N__4735));
    LocalMux I__500 (
            .O(N__4738),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    LocalMux I__499 (
            .O(N__4735),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ));
    IoInMux I__498 (
            .O(N__4730),
            .I(N__4727));
    LocalMux I__497 (
            .O(N__4727),
            .I(N__4724));
    IoSpan4Mux I__496 (
            .O(N__4724),
            .I(N__4721));
    IoSpan4Mux I__495 (
            .O(N__4721),
            .I(N__4718));
    Span4Mux_s2_v I__494 (
            .O(N__4718),
            .I(N__4714));
    InMux I__493 (
            .O(N__4717),
            .I(N__4711));
    Sp12to4 I__492 (
            .O(N__4714),
            .I(N__4708));
    LocalMux I__491 (
            .O(N__4711),
            .I(N__4705));
    Span12Mux_s8_v I__490 (
            .O(N__4708),
            .I(N__4702));
    Span4Mux_h I__489 (
            .O(N__4705),
            .I(N__4699));
    Span12Mux_v I__488 (
            .O(N__4702),
            .I(N__4694));
    Sp12to4 I__487 (
            .O(N__4699),
            .I(N__4694));
    Odrv12 I__486 (
            .O(N__4694),
            .I(A_c_10));
    CascadeMux I__485 (
            .O(N__4691),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ));
    InMux I__484 (
            .O(N__4688),
            .I(N__4685));
    LocalMux I__483 (
            .O(N__4685),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ));
    InMux I__482 (
            .O(N__4682),
            .I(N__4679));
    LocalMux I__481 (
            .O(N__4679),
            .I(N__4676));
    Odrv4 I__480 (
            .O(N__4676),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ));
    IoInMux I__479 (
            .O(N__4673),
            .I(N__4670));
    LocalMux I__478 (
            .O(N__4670),
            .I(N__4667));
    IoSpan4Mux I__477 (
            .O(N__4667),
            .I(N__4664));
    Sp12to4 I__476 (
            .O(N__4664),
            .I(N__4661));
    Span12Mux_s7_h I__475 (
            .O(N__4661),
            .I(N__4658));
    Span12Mux_h I__474 (
            .O(N__4658),
            .I(N__4655));
    Odrv12 I__473 (
            .O(N__4655),
            .I(CMA_c_7));
    IoInMux I__472 (
            .O(N__4652),
            .I(N__4649));
    LocalMux I__471 (
            .O(N__4649),
            .I(N__4646));
    IoSpan4Mux I__470 (
            .O(N__4646),
            .I(N__4643));
    Sp12to4 I__469 (
            .O(N__4643),
            .I(N__4640));
    Span12Mux_s7_h I__468 (
            .O(N__4640),
            .I(N__4637));
    Span12Mux_h I__467 (
            .O(N__4637),
            .I(N__4634));
    Odrv12 I__466 (
            .O(N__4634),
            .I(CMA_c_8));
    InMux I__465 (
            .O(N__4631),
            .I(N__4628));
    LocalMux I__464 (
            .O(N__4628),
            .I(\U712_CHIP_RAM.REFRESH5lto0 ));
    InMux I__463 (
            .O(N__4625),
            .I(bfn_9_5_0_));
    InMux I__462 (
            .O(N__4622),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ));
    InMux I__461 (
            .O(N__4619),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ));
    InMux I__460 (
            .O(N__4616),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ));
    InMux I__459 (
            .O(N__4613),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ));
    InMux I__458 (
            .O(N__4610),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ));
    InMux I__457 (
            .O(N__4607),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ));
    InMux I__456 (
            .O(N__4604),
            .I(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ));
    ClkMux I__455 (
            .O(N__4601),
            .I(N__4586));
    ClkMux I__454 (
            .O(N__4600),
            .I(N__4586));
    ClkMux I__453 (
            .O(N__4599),
            .I(N__4586));
    ClkMux I__452 (
            .O(N__4598),
            .I(N__4586));
    ClkMux I__451 (
            .O(N__4597),
            .I(N__4586));
    GlobalMux I__450 (
            .O(N__4586),
            .I(N__4583));
    gio2CtrlBuf I__449 (
            .O(N__4583),
            .I(C1_c_g));
    InMux I__448 (
            .O(N__4580),
            .I(N__4576));
    InMux I__447 (
            .O(N__4579),
            .I(N__4573));
    LocalMux I__446 (
            .O(N__4576),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    LocalMux I__445 (
            .O(N__4573),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ));
    InMux I__444 (
            .O(N__4568),
            .I(N__4564));
    InMux I__443 (
            .O(N__4567),
            .I(N__4561));
    LocalMux I__442 (
            .O(N__4564),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    LocalMux I__441 (
            .O(N__4561),
            .I(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ));
    IoInMux I__440 (
            .O(N__4556),
            .I(N__4553));
    LocalMux I__439 (
            .O(N__4553),
            .I(N__4550));
    Span4Mux_s0_v I__438 (
            .O(N__4550),
            .I(N__4547));
    Span4Mux_v I__437 (
            .O(N__4547),
            .I(N__4544));
    Span4Mux_v I__436 (
            .O(N__4544),
            .I(N__4541));
    Span4Mux_v I__435 (
            .O(N__4541),
            .I(N__4538));
    Odrv4 I__434 (
            .O(N__4538),
            .I(CMA_c_1));
    InMux I__433 (
            .O(N__4535),
            .I(N__4532));
    LocalMux I__432 (
            .O(N__4532),
            .I(\U712_CHIP_RAM.N_340 ));
    IoInMux I__431 (
            .O(N__4529),
            .I(N__4526));
    LocalMux I__430 (
            .O(N__4526),
            .I(N__4523));
    IoSpan4Mux I__429 (
            .O(N__4523),
            .I(N__4520));
    Span4Mux_s3_h I__428 (
            .O(N__4520),
            .I(N__4517));
    Sp12to4 I__427 (
            .O(N__4517),
            .I(N__4514));
    Span12Mux_s8_h I__426 (
            .O(N__4514),
            .I(N__4511));
    Span12Mux_h I__425 (
            .O(N__4511),
            .I(N__4508));
    Odrv12 I__424 (
            .O(N__4508),
            .I(CMA_c_5));
    InMux I__423 (
            .O(N__4505),
            .I(N__4502));
    LocalMux I__422 (
            .O(N__4502),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ));
    CascadeMux I__421 (
            .O(N__4499),
            .I(\U712_CHIP_RAM.N_297_cascade_ ));
    InMux I__420 (
            .O(N__4496),
            .I(N__4493));
    LocalMux I__419 (
            .O(N__4493),
            .I(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ));
    CascadeMux I__418 (
            .O(N__4490),
            .I(\U712_CHIP_RAM.N_196_cascade_ ));
    IoInMux I__417 (
            .O(N__4487),
            .I(N__4483));
    IoInMux I__416 (
            .O(N__4486),
            .I(N__4480));
    LocalMux I__415 (
            .O(N__4483),
            .I(N__4477));
    LocalMux I__414 (
            .O(N__4480),
            .I(N__4474));
    Span4Mux_s2_v I__413 (
            .O(N__4477),
            .I(N__4471));
    IoSpan4Mux I__412 (
            .O(N__4474),
            .I(N__4468));
    Span4Mux_h I__411 (
            .O(N__4471),
            .I(N__4465));
    Span4Mux_s2_v I__410 (
            .O(N__4468),
            .I(N__4462));
    Sp12to4 I__409 (
            .O(N__4465),
            .I(N__4458));
    Span4Mux_h I__408 (
            .O(N__4462),
            .I(N__4455));
    IoInMux I__407 (
            .O(N__4461),
            .I(N__4452));
    Span12Mux_h I__406 (
            .O(N__4458),
            .I(N__4447));
    Sp12to4 I__405 (
            .O(N__4455),
            .I(N__4447));
    LocalMux I__404 (
            .O(N__4452),
            .I(N__4444));
    Span12Mux_v I__403 (
            .O(N__4447),
            .I(N__4438));
    Span12Mux_s11_h I__402 (
            .O(N__4444),
            .I(N__4438));
    InMux I__401 (
            .O(N__4443),
            .I(N__4435));
    Odrv12 I__400 (
            .O(N__4438),
            .I(TACK_EN));
    LocalMux I__399 (
            .O(N__4435),
            .I(TACK_EN));
    IoInMux I__398 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__397 (
            .O(N__4427),
            .I(N__4424));
    Span12Mux_s6_v I__396 (
            .O(N__4424),
            .I(N__4421));
    Odrv12 I__395 (
            .O(N__4421),
            .I(CLK80_PLL_i_i));
    IoInMux I__394 (
            .O(N__4418),
            .I(N__4415));
    LocalMux I__393 (
            .O(N__4415),
            .I(N__4412));
    Span4Mux_s3_h I__392 (
            .O(N__4412),
            .I(N__4409));
    Odrv4 I__391 (
            .O(N__4409),
            .I(DBRn_c_i_0));
    IoInMux I__390 (
            .O(N__4406),
            .I(N__4403));
    LocalMux I__389 (
            .O(N__4403),
            .I(N__4400));
    Span12Mux_s3_v I__388 (
            .O(N__4400),
            .I(N__4397));
    Odrv12 I__387 (
            .O(N__4397),
            .I(VBENn_c));
    InMux I__386 (
            .O(N__4394),
            .I(N__4391));
    LocalMux I__385 (
            .O(N__4391),
            .I(N__4388));
    Span4Mux_h I__384 (
            .O(N__4388),
            .I(N__4385));
    Sp12to4 I__383 (
            .O(N__4385),
            .I(N__4382));
    Span12Mux_v I__382 (
            .O(N__4382),
            .I(N__4379));
    Odrv12 I__381 (
            .O(N__4379),
            .I(A_c_14));
    IoInMux I__380 (
            .O(N__4376),
            .I(N__4373));
    LocalMux I__379 (
            .O(N__4373),
            .I(N__4370));
    IoSpan4Mux I__378 (
            .O(N__4370),
            .I(N__4367));
    Span4Mux_s2_v I__377 (
            .O(N__4367),
            .I(N__4364));
    Sp12to4 I__376 (
            .O(N__4364),
            .I(N__4361));
    Span12Mux_v I__375 (
            .O(N__4361),
            .I(N__4358));
    Odrv12 I__374 (
            .O(N__4358),
            .I(CLK40_IN_c));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .I(N__4600));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .I(N__4597));
    INV \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C  (
            .O(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .I(N__4598));
    INV \INVU712_CHIP_RAM.DMA_A1_nesrC  (
            .O(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .I(N__4599));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_10_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_12_0_));
    ICE_GB C1_ibuf_RNIPA2A (
            .USERSIGNALTOGLOBALBUFFER(N__5434),
            .GLOBALBUFFEROUTPUT(C1_c_g));
    ICE_GB RESETn_ibuf_RNIM9SF_0 (
            .USERSIGNALTOGLOBALBUFFER(N__8636),
            .GLOBALBUFFEROUTPUT(RESETn_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    ICE_GB DBRn_c_i_0_g_gb (
            .USERSIGNALTOGLOBALBUFFER(N__4418),
            .GLOBALBUFFEROUTPUT(DBRn_c_i_0_g));
    ICE_GB C3_ibuf_RNIRKME (
            .USERSIGNALTOGLOBALBUFFER(N__5105),
            .GLOBALBUFFEROUTPUT(C3_c_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam CLKRAM_obuf_RNO_LC_2_1_6.C_ON=1'b0;
    defparam CLKRAM_obuf_RNO_LC_2_1_6.SEQ_MODE=4'b0000;
    defparam CLKRAM_obuf_RNO_LC_2_1_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 CLKRAM_obuf_RNO_LC_2_1_6 (
            .in0(N__10274),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK80_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_3_11_2  (
            .in0(_gnd_net_),
            .in1(N__10736),
            .in2(_gnd_net_),
            .in3(N__8725),
            .lcout(DBRn_c_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.C_ON=1'b0;
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.SEQ_MODE=4'b0000;
    defparam DBRn_ibuf_RNIBAB_LC_6_14_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBRn_ibuf_RNIBAB_LC_6_14_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5188),
            .lcout(DBRn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_4 .C_ON=1'b0;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_BUFFERS.un1_VBENn_0_a2_LC_8_6_4  (
            .in0(N__10042),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10126),
            .lcout(VBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_6_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_8_6_7  (
            .in0(N__4394),
            .in1(N__10041),
            .in2(_gnd_net_),
            .in3(N__9032),
            .lcout(\U712_CHIP_RAM.N_340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_8_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_1_LC_8_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_1_LC_8_7_5  (
            .in0(N__4505),
            .in1(N__4496),
            .in2(_gnd_net_),
            .in3(N__4688),
            .lcout(CMA_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10246),
            .ce(N__11217),
            .sr(N__10700));
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_8_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_5_LC_8_7_6 .LUT_INIT=16'b1000111110000101;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_5_LC_8_7_6  (
            .in0(N__8549),
            .in1(N__4535),
            .in2(N__9225),
            .in3(N__5537),
            .lcout(CMA_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10246),
            .ce(N__11217),
            .sr(N__10700));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_8_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_8_8_0 .LUT_INIT=16'b1110111100001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_8_8_0  (
            .in0(N__10050),
            .in1(N__8768),
            .in2(N__9226),
            .in3(N__8548),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_8_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_8_8_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__5668),
            .in2(_gnd_net_),
            .in3(N__6889),
            .lcout(\U712_CHIP_RAM.N_297 ),
            .ltout(\U712_CHIP_RAM.N_297_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_8_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_8_8_2 .LUT_INIT=16'b0100000000001111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_8_8_2  (
            .in0(N__10051),
            .in1(N__8767),
            .in2(N__4499),
            .in3(N__9214),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_9_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_9_0  (
            .in0(N__4883),
            .in1(N__7599),
            .in2(N__7703),
            .in3(N__4859),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_TACK_LC_8_9_1 .LUT_INIT=16'b1010110010101111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_LC_8_9_1  (
            .in0(N__5871),
            .in1(N__5738),
            .in2(N__4490),
            .in3(N__8139),
            .lcout(CPU_TACKm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10253),
            .ce(),
            .sr(N__10687));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_8_9_4  (
            .in0(N__7468),
            .in1(N__7598),
            .in2(N__8051),
            .in3(N__7329),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_9_7 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_8_9_7  (
            .in0(N__4877),
            .in1(N__5602),
            .in2(_gnd_net_),
            .in3(N__6479),
            .lcout(\U712_CHIP_RAM.N_202 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_LC_8_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_8_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_EN_LC_8_13_0 .LUT_INIT=16'b0100010011111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_LC_8_13_0  (
            .in0(N__5155),
            .in1(N__4443),
            .in2(_gnd_net_),
            .in3(N__5282),
            .lcout(TACK_EN),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10267),
            .ce(),
            .sr(N__10667));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_5_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_5_0 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__4631),
            .in2(_gnd_net_),
            .in3(N__4625),
            .lcout(\U712_CHIP_RAM.REFRESH5lto0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_5_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__4568),
            .in2(_gnd_net_),
            .in3(N__4622),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_5_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_5_2 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__4787),
            .in2(_gnd_net_),
            .in3(N__4619),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_5_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_5_3 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__4580),
            .in2(_gnd_net_),
            .in3(N__4616),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_5_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_5_4 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__4801),
            .in2(_gnd_net_),
            .in3(N__4613),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_5_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_5_5 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__4742),
            .in2(_gnd_net_),
            .in3(N__4610),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_5_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_5_6 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__4754),
            .in2(_gnd_net_),
            .in3(N__4607),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.REFRESH_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.REFRESH_COUNTER_cry_6 ),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_5_7 .SEQ_MODE=4'b1010;
    defparam \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_5_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__4852),
            .in2(_gnd_net_),
            .in3(N__4604),
            .lcout(\U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4601),
            .ce(),
            .sr(N__5468));
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_6_0 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_0_LC_9_6_0  (
            .in0(N__4579),
            .in1(N__4567),
            .in2(N__4802),
            .in3(N__4786),
            .lcout(\U712_CHIP_RAM.REFRESH5lt7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_9_6_2  (
            .in0(N__4775),
            .in1(N__7097),
            .in2(_gnd_net_),
            .in3(N__9167),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_9_6_3  (
            .in0(N__9169),
            .in1(N__10029),
            .in2(N__4757),
            .in3(N__8741),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_6_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CHIP_RAM.REFRESH_RNO_1_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__4753),
            .in2(_gnd_net_),
            .in3(N__4741),
            .lcout(\U712_CHIP_RAM.REFRESH5lto7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_9_6_6  (
            .in0(N__4717),
            .in1(N__7214),
            .in2(_gnd_net_),
            .in3(N__9166),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_6_7 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_9_6_7  (
            .in0(N__9168),
            .in1(N__10028),
            .in2(N__4691),
            .in3(N__8822),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_9_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_7_LC_9_7_3 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_7_LC_9_7_3  (
            .in0(N__8550),
            .in1(N__8831),
            .in2(N__8521),
            .in3(N__4682),
            .lcout(CMA_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10240),
            .ce(N__11195),
            .sr(N__10695));
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_8_LC_9_7_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_8_LC_9_7_6  (
            .in0(N__8551),
            .in1(N__8753),
            .in2(N__8522),
            .in3(N__5543),
            .lcout(CMA_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10240),
            .ce(N__11195),
            .sr(N__10695));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_7_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_LC_9_7_7  (
            .in0(N__5667),
            .in1(N__9137),
            .in2(N__6897),
            .in3(N__5491),
            .lcout(\U712_CHIP_RAM.REFRESH_RST ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_1 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_0_LC_9_8_1  (
            .in0(N__4910),
            .in1(N__5523),
            .in2(N__6901),
            .in3(N__5637),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10247),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_8_2 .LUT_INIT=16'b0000110011101010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_2_LC_9_8_2  (
            .in0(N__8038),
            .in1(N__7589),
            .in2(N__8153),
            .in3(N__7323),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_95_i_a2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_3 .LUT_INIT=16'b1111000011100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_3_LC_9_8_3  (
            .in0(N__5588),
            .in1(N__5524),
            .in2(N__5509),
            .in3(N__5638),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10247),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_8_4 .LUT_INIT=16'b0100010001000101;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIVA2D1_LC_9_8_4  (
            .in0(N__6967),
            .in1(N__5063),
            .in2(N__4820),
            .in3(N__4934),
            .lcout(\U712_CHIP_RAM.N_556 ),
            .ltout(\U712_CHIP_RAM.N_556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_8_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_0_2_LC_9_8_5  (
            .in0(N__10567),
            .in1(N__8039),
            .in2(N__4871),
            .in3(N__6455),
            .lcout(\U712_CHIP_RAM.N_388 ),
            .ltout(\U712_CHIP_RAM.N_388_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6 .LUT_INIT=16'b1111111000000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_2_LC_9_8_6  (
            .in0(N__5636),
            .in1(N__4868),
            .in2(N__4862),
            .in3(N__5671),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10247),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_7 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_9_8_7  (
            .in0(N__7588),
            .in1(N__4819),
            .in2(N__8050),
            .in3(N__6968),
            .lcout(\U712_CHIP_RAM.N_445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_0 .LUT_INIT=16'b1001010110010111;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_9_9_0  (
            .in0(N__8150),
            .in1(N__7897),
            .in2(N__7333),
            .in3(N__7469),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNIIICT_LC_9_9_1  (
            .in0(N__4815),
            .in1(N__5059),
            .in2(_gnd_net_),
            .in3(N__4932),
            .lcout(\U712_CHIP_RAM.N_551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.REFRESH_LC_9_9_2 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \U712_CHIP_RAM.REFRESH_LC_9_9_2  (
            .in0(N__4853),
            .in1(N__4838),
            .in2(N__10568),
            .in3(N__4829),
            .lcout(\U712_CHIP_RAM.REFRESHZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10250),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMM5O1_3_LC_9_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMM5O1_3_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIMM5O1_3_LC_9_9_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIMM5O1_3_LC_9_9_3  (
            .in0(N__7587),
            .in1(N__7324),
            .in2(N__7905),
            .in3(N__8149),
            .lcout(\U712_CHIP_RAM.N_303 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4 .LUT_INIT=16'b1100110000001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_LC_9_9_4  (
            .in0(N__6984),
            .in1(N__10562),
            .in2(N__11174),
            .in3(N__4904),
            .lcout(\U712_CHIP_RAM.DMA_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10250),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(N__10052),
            .in2(_gnd_net_),
            .in3(N__4933),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_417_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6 .LUT_INIT=16'b1111000100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_START_LC_9_9_6  (
            .in0(N__4952),
            .in1(N__5018),
            .in2(N__4937),
            .in3(N__10561),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10250),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_9_7 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_9_9_7  (
            .in0(N__10563),
            .in1(N__6278),
            .in2(N__4919),
            .in3(N__7699),
            .lcout(\U712_CHIP_RAM.N_206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_9_10_0  (
            .in0(N__4898),
            .in1(N__4891),
            .in2(_gnd_net_),
            .in3(N__5941),
            .lcout(\U712_CHIP_RAM.N_457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_10_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_5_LC_9_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_5_LC_9_10_2  (
            .in0(N__10560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4892),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10254),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_4_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__10559),
            .in2(_gnd_net_),
            .in3(N__7715),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10254),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_10_6 .LUT_INIT=16'b1100110011011101;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_9_10_6  (
            .in0(N__10049),
            .in1(N__5783),
            .in2(_gnd_net_),
            .in3(N__7385),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_8_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_7 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_LC_9_10_7  (
            .in0(N__5942),
            .in1(N__5847),
            .in2(N__5753),
            .in3(N__10558),
            .lcout(\U712_CHIP_RAM.RAM_CYCLE_DISABLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10254),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_11_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.LATCH_CLK_LC_9_11_7 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_LC_9_11_7  (
            .in0(N__11168),
            .in1(N__5765),
            .in2(N__7334),
            .in3(N__5029),
            .lcout(LATCH_CLK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10257),
            .ce(),
            .sr(N__10670));
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_1_LC_9_12_0  (
            .in0(N__10549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6629),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10262),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_7 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_START_LC_9_12_7 .LUT_INIT=16'b1100110000000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_LC_9_12_7  (
            .in0(N__5011),
            .in1(N__10550),
            .in2(N__4985),
            .in3(N__4961),
            .lcout(\U712_REG_SM.REG_CYCLE_STARTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10262),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_3_LC_9_13_0  (
            .in0(N__5276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10553),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10265),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_13_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_START_RNO_0_LC_9_13_1  (
            .in0(N__5446),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6093),
            .lcout(\U712_REG_SM.N_414 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_13_2 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_13_2 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_9_13_2  (
            .in0(N__5116),
            .in1(N__5141),
            .in2(N__5885),
            .in3(N__6542),
            .lcout(),
            .ltout(\U712_CYCLE_TERM.N_452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_3 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_3 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_3 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_1_LC_9_13_3  (
            .in0(N__10551),
            .in1(N__9528),
            .in2(N__4955),
            .in3(N__5117),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10265),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_4 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_4 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_2_LC_9_13_4  (
            .in0(N__9527),
            .in1(N__10552),
            .in2(_gnd_net_),
            .in3(N__5142),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10265),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_13_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_13_5 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \U712_CYCLE_TERM.TACK_EN_RNO_0_LC_9_13_5  (
            .in0(N__6541),
            .in1(N__5881),
            .in2(_gnd_net_),
            .in3(N__5115),
            .lcout(\U712_CYCLE_TERM.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_4_LC_9_13_6  (
            .in0(N__5266),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10554),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10265),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_13_7 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_13_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_1_0_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__5265),
            .in2(_gnd_net_),
            .in3(N__5275),
            .lcout(\U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_0 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_0 .LUT_INIT=16'b1111111111000100;
    LogicCell40 \U712_CYCLE_TERM.TACK_OUTn_LC_9_14_0  (
            .in0(N__5144),
            .in1(N__5205),
            .in2(N__9530),
            .in3(N__5267),
            .lcout(TACK_OUTn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_1_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_1_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5399),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam DBR_SYNC_0_LC_9_14_3.C_ON=1'b0;
    defparam DBR_SYNC_0_LC_9_14_3.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_0_LC_9_14_3.LUT_INIT=16'b1010101010101010;
    LogicCell40 DBR_SYNC_0_LC_9_14_3 (
            .in0(N__5192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(DBR_SYNCZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam DBR_SYNC_1_LC_9_14_4.C_ON=1'b0;
    defparam DBR_SYNC_1_LC_9_14_4.SEQ_MODE=4'b1001;
    defparam DBR_SYNC_1_LC_9_14_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 DBR_SYNC_1_LC_9_14_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5162),
            .lcout(DBR_SYNCZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_5 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_5 .LUT_INIT=16'b0011001000100010;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_0_LC_9_14_5  (
            .in0(N__5156),
            .in1(N__5143),
            .in2(N__5126),
            .in3(N__5855),
            .lcout(\U712_CYCLE_TERM.TACK_STATEZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_0_LC_9_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_REG_SM.C3_SYNC_0_LC_9_14_6  (
            .in0(N__5092),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam \U712_REG_SM.START_RST_LC_9_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.START_RST_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.START_RST_LC_9_14_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \U712_REG_SM.START_RST_LC_9_14_7  (
            .in0(N__6618),
            .in1(N__5447),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(\U712_REG_SM.START_RSTZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10268),
            .ce(),
            .sr(N__10665));
    defparam \U712_REG_SM.REGENn_LC_9_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_LC_9_15_1 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.REGENn_LC_9_15_1 .LUT_INIT=16'b1010011010100010;
    LogicCell40 \U712_REG_SM.REGENn_LC_9_15_1  (
            .in0(N__6124),
            .in1(N__6107),
            .in2(N__9365),
            .in3(N__6737),
            .lcout(REGENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10269),
            .ce(),
            .sr(N__10664));
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_15_2 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C1_SYNC_0_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C1_SYNC_0_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5435),
            .lcout(\U712_REG_SM.C1_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10269),
            .ce(),
            .sr(N__10664));
    defparam \U712_CHIP_RAM.CRCSn_LC_10_1_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CRCSn_LC_10_1_3 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CRCSn_LC_10_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CRCSn_LC_10_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5510),
            .lcout(CRCSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10225),
            .ce(),
            .sr(N__10707));
    defparam \U712_CHIP_RAM.RASn_LC_10_4_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RASn_LC_10_4_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.RASn_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.RASn_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5678),
            .lcout(RASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10229),
            .ce(),
            .sr(N__10703));
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_10_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_10_5_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_0_LC_10_5_0 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_0_LC_10_5_0  (
            .in0(N__8511),
            .in1(N__8569),
            .in2(N__5576),
            .in3(N__8885),
            .lcout(CMA_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(N__11207),
            .sr(N__10701));
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_5_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_10_LC_10_5_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_10_LC_10_5_6  (
            .in0(N__9224),
            .in1(N__5508),
            .in2(_gnd_net_),
            .in3(N__8570),
            .lcout(CMA_c_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(N__11207),
            .sr(N__10701));
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_10_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_2_LC_10_5_7 .LUT_INIT=16'b1010001010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_2_LC_10_5_7  (
            .in0(N__8571),
            .in1(N__8512),
            .in2(N__8984),
            .in3(N__6266),
            .lcout(CMA_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10232),
            .ce(N__11207),
            .sr(N__10701));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_6_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_10_6_0  (
            .in0(N__6752),
            .in1(N__5317),
            .in2(_gnd_net_),
            .in3(N__9162),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_1 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_10_6_1  (
            .in0(N__9164),
            .in1(N__10000),
            .in2(N__5579),
            .in3(N__8423),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_6_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_6_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_8_LC_10_6_2  (
            .in0(N__5567),
            .in1(N__6193),
            .in2(_gnd_net_),
            .in3(N__9163),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_6_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_6_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_8_LC_10_6_3  (
            .in0(N__9165),
            .in1(N__10001),
            .in2(N__5546),
            .in3(N__8702),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_6_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_10_6_5  (
            .in0(N__7154),
            .in1(N__9999),
            .in2(_gnd_net_),
            .in3(N__8792),
            .lcout(\U712_CHIP_RAM.N_346 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_0 .LUT_INIT=16'b1010101010111000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_1_LC_10_7_0  (
            .in0(N__9152),
            .in1(N__5639),
            .in2(N__5612),
            .in3(N__5525),
            .lcout(\U712_CHIP_RAM.SDRAM_CMDZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10238),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_7_1 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNI32HB1_3_LC_10_7_1  (
            .in0(N__5669),
            .in1(N__9150),
            .in2(N__5504),
            .in3(N__5464),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_CMA25_0_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_7_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNIPBDR1_3_LC_10_7_2  (
            .in0(N__10734),
            .in1(_gnd_net_),
            .in2(N__5450),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_CMA25_0_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_7_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNO_0_LC_10_7_4  (
            .in0(N__10735),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7485),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_7_5 .LUT_INIT=16'b1101110001010000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_1_LC_10_7_5  (
            .in0(N__6985),
            .in1(N__7420),
            .in2(N__7489),
            .in3(N__7628),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_7_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_7_6 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNO_0_LC_10_7_6  (
            .in0(N__10733),
            .in1(_gnd_net_),
            .in2(N__5681),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_10_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_10_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_10_7_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_10_7_7 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_9_LC_10_7_7  (
            .in0(N__5670),
            .in1(N__9151),
            .in2(_gnd_net_),
            .in3(N__6890),
            .lcout(\U712_CHIP_RAM.CMA_5_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_8_0 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIEVI78_3_LC_10_8_0  (
            .in0(N__10548),
            .in1(N__7906),
            .in2(N__6338),
            .in3(N__6500),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_8_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_10_8_1  (
            .in0(N__6325),
            .in1(N__6485),
            .in2(N__5621),
            .in3(N__6474),
            .lcout(\U712_CHIP_RAM.N_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_8_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_1_3_LC_10_8_2  (
            .in0(N__7576),
            .in1(_gnd_net_),
            .in2(N__8152),
            .in3(N__8022),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_443_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_3  (
            .in0(N__6326),
            .in1(N__5603),
            .in2(N__5591),
            .in3(N__6475),
            .lcout(\U712_CHIP_RAM.N_204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_0_LC_10_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_0_LC_10_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_0_LC_10_8_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_0_LC_10_8_4  (
            .in0(_gnd_net_),
            .in1(N__7467),
            .in2(_gnd_net_),
            .in3(N__8021),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIVSQ24_LC_10_8_5  (
            .in0(N__7675),
            .in1(N__6363),
            .in2(N__6312),
            .in3(N__7575),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_10_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_10_8_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI05TJ3_LC_10_8_6  (
            .in0(N__7574),
            .in1(N__6301),
            .in2(N__8151),
            .in3(N__7676),
            .lcout(\U712_CHIP_RAM.N_463 ),
            .ltout(\U712_CHIP_RAM.N_463_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_8_7 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNIU7TF5_LC_10_8_7  (
            .in0(N__8020),
            .in1(N__6966),
            .in2(N__5582),
            .in3(N__6253),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_10_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_10_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_10_9_0 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_1_LC_10_9_0  (
            .in0(N__7590),
            .in1(N__6509),
            .in2(N__7349),
            .in3(N__7684),
            .lcout(),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_10_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_10_9_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_0_LC_10_9_1  (
            .in0(N__10730),
            .in1(_gnd_net_),
            .in2(N__5741),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI9UML3_LC_10_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI9UML3_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI9UML3_LC_10_9_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI9UML3_LC_10_9_2  (
            .in0(N__11131),
            .in1(N__7376),
            .in2(_gnd_net_),
            .in3(N__6499),
            .lcout(\U712_CHIP_RAM.N_418 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_9_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_10_9_3  (
            .in0(N__7685),
            .in1(N__10059),
            .in2(N__6316),
            .in3(N__8043),
            .lcout(\U712_CHIP_RAM.N_439 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_4 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_10_9_4  (
            .in0(N__7591),
            .in1(N__6347),
            .in2(_gnd_net_),
            .in3(N__10545),
            .lcout(\U712_CHIP_RAM.SDRAM_CONFIGUREDZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10248),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_9_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_START_RNICLGI4_LC_10_9_5  (
            .in0(N__6986),
            .in1(N__8042),
            .in2(_gnd_net_),
            .in3(N__6454),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1 ),
            .ltout(\U712_CHIP_RAM.WRITE_CYCLE_0_sqmuxa_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_9_6 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNIMAOKC_LC_10_9_6  (
            .in0(N__5729),
            .in1(N__5776),
            .in2(N__5723),
            .in3(N__7623),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0 ),
            .ltout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_9_7 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_10_9_7  (
            .in0(N__10731),
            .in1(_gnd_net_),
            .in2(N__5720),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_10_0 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CLK_EN_ess_LC_10_10_0 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_LC_10_10_0  (
            .in0(N__6368),
            .in1(_gnd_net_),
            .in2(N__7907),
            .in3(N__7328),
            .lcout(CLK_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10251),
            .ce(N__5693),
            .sr(N__10671));
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_10_1 .LUT_INIT=16'b1110111000110011;
    LogicCell40 \U712_CHIP_RAM.CPU_TACK_RNO_4_LC_10_10_1  (
            .in0(N__7466),
            .in1(N__8041),
            .in2(_gnd_net_),
            .in3(N__7901),
            .lcout(\U712_CHIP_RAM.N_360 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_10_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_10_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \U712_CHIP_RAM.LATCH_CLK_RNO_0_LC_10_10_3  (
            .in0(N__7421),
            .in1(N__5777),
            .in2(_gnd_net_),
            .in3(N__7627),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_10_11_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_10_11_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_2_LC_10_11_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_2_LC_10_11_0  (
            .in0(N__5841),
            .in1(N__10412),
            .in2(N__5990),
            .in3(N__5937),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10255),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_11_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_11_2 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_11_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_3_LC_10_11_2  (
            .in0(N__6575),
            .in1(N__6156),
            .in2(N__5848),
            .in3(N__8299),
            .lcout(),
            .ltout(\U712_REG_SM.N_400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_11_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_3_LC_10_11_3 .LUT_INIT=16'b0000101000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_3_LC_10_11_3  (
            .in0(N__10413),
            .in1(N__8303),
            .in2(N__5759),
            .in3(N__9364),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10255),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_11_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_11_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_1_LC_10_11_6  (
            .in0(N__5971),
            .in1(N__6001),
            .in2(N__5900),
            .in3(N__5936),
            .lcout(),
            .ltout(\U712_CHIP_RAM.RAM_CYCLE_DISABLE_6_iv_i_a2_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_11_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_11_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_11_7 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \U712_CHIP_RAM.RAM_CYCLE_DISABLE_RNO_0_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(N__5954),
            .in2(N__5756),
            .in3(N__5837),
            .lcout(\U712_CHIP_RAM.N_405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_10_12_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_10_12_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_0_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(N__5896),
            .in2(N__5798),
            .in3(N__5797),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_10_12_0_),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_10_12_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_10_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_10_12_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_1_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(N__5953),
            .in2(_gnd_net_),
            .in3(N__5744),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_10_12_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_10_12_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_2_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(N__6002),
            .in2(_gnd_net_),
            .in3(N__5981),
            .lcout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.un1_CAS_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_10_12_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_10_12_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_RNO_0_3_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(N__5972),
            .in2(_gnd_net_),
            .in3(N__5978),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CAS_COUNTER_RNO_0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_10_12_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_3_LC_10_12_4 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_3_LC_10_12_4  (
            .in0(N__5939),
            .in1(N__10489),
            .in2(N__5975),
            .in3(N__5846),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10258),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_10_12_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_1_LC_10_12_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_1_LC_10_12_5  (
            .in0(N__10488),
            .in1(N__5940),
            .in2(N__5849),
            .in3(N__5960),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10258),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_10_12_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_10_12_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_COUNTER_0_LC_10_12_6 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_CHIP_RAM.CAS_COUNTER_0_LC_10_12_6  (
            .in0(N__5938),
            .in1(N__5845),
            .in2(N__5909),
            .in3(N__10487),
            .lcout(\U712_CHIP_RAM.CAS_COUNTERZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10258),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_13_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_13_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNIH4AH_1_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(N__8280),
            .in2(_gnd_net_),
            .in3(N__5819),
            .lcout(\U712_REG_SM.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_13_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3OIA1_0_LC_10_13_4  (
            .in0(N__6728),
            .in1(N__6094),
            .in2(N__8297),
            .in3(N__9326),
            .lcout(\U712_REG_SM.STATE_COUNT_0_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_6 .C_ON=1'b0;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_10_13_6  (
            .in0(N__6531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5880),
            .lcout(\U712_CYCLE_TERM.TACK_EN6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam DBR_SYNC_RNITKK4_1_LC_10_13_7.C_ON=1'b0;
    defparam DBR_SYNC_RNITKK4_1_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam DBR_SYNC_RNITKK4_1_LC_10_13_7.LUT_INIT=16'b0000000011111111;
    LogicCell40 DBR_SYNC_RNITKK4_1_LC_10_13_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5818),
            .lcout(DBR_SYNC_i_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_10_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_10_14_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__9325),
            .in2(_gnd_net_),
            .in3(N__8275),
            .lcout(\U712_REG_SM.N_307 ),
            .ltout(\U712_REG_SM.N_307_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_14_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_1_LC_10_14_1  (
            .in0(N__8220),
            .in1(N__10112),
            .in2(N__6161),
            .in3(N__6077),
            .lcout(\U712_REG_SM.REG_CYCLE_5_iv_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_10_14_3 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_10_14_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNIJUGT_3_LC_10_14_3  (
            .in0(N__8276),
            .in1(N__9327),
            .in2(_gnd_net_),
            .in3(N__6158),
            .lcout(\U712_REG_SM.N_553 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_0_LC_10_14_4  (
            .in0(N__6076),
            .in1(N__6157),
            .in2(_gnd_net_),
            .in3(N__8221),
            .lcout(\U712_REG_SM.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REGENn_RNO_0_LC_10_15_1 .LUT_INIT=16'b0000110001010000;
    LogicCell40 \U712_REG_SM.REGENn_RNO_0_LC_10_15_1  (
            .in0(N__6100),
            .in1(N__8338),
            .in2(N__8298),
            .in3(N__6123),
            .lcout(\U712_REG_SM.REGENn_e_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_15_7 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_15_7 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_0_LC_10_15_7  (
            .in0(N__6101),
            .in1(N__8284),
            .in2(N__9352),
            .in3(N__6729),
            .lcout(\U712_REG_SM.STATE_COUNTsr_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_16_6 .C_ON=1'b0;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_16_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.WRITE_CYCLE_LC_10_16_6 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_REG_SM.WRITE_CYCLE_LC_10_16_6  (
            .in0(N__9808),
            .in1(N__6075),
            .in2(_gnd_net_),
            .in3(N__6620),
            .lcout(\U712_REG_SM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10270),
            .ce(),
            .sr(N__10661));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_5_2 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_11_5_2  (
            .in0(N__6059),
            .in1(N__7070),
            .in2(N__9209),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_4 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_11_5_4  (
            .in0(N__6037),
            .in1(N__7181),
            .in2(N__9210),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_5 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_11_5_5  (
            .in0(N__9220),
            .in1(N__9993),
            .in2(N__6269),
            .in3(N__9668),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_5_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEA_LC_11_5_7  (
            .in0(_gnd_net_),
            .in1(N__9992),
            .in2(_gnd_net_),
            .in3(N__9173),
            .lcout(\U712_CHIP_RAM.CPU_CYCLE_esr_RNIHMEAZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_6_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_CHIP_RAM.CPU_CYCLE_esr_LC_11_6_0  (
            .in0(N__6997),
            .in1(N__6179),
            .in2(_gnd_net_),
            .in3(N__6260),
            .lcout(CPU_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10233),
            .ce(N__6242),
            .sr(N__10688));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_0_LC_11_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_0_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_0_LC_11_7_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_0_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__6229),
            .in2(_gnd_net_),
            .in3(N__10732),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_11_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_11_7_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_1_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__7980),
            .in2(_gnd_net_),
            .in3(N__8124),
            .lcout(\U712_CHIP_RAM.N_302 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_7_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_8_LC_11_7_3  (
            .in0(N__6230),
            .in1(N__6215),
            .in2(N__10997),
            .in3(N__6194),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10236),
            .ce(),
            .sr(N__10680));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_7_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI5KG83_1_LC_11_7_4  (
            .in0(N__7692),
            .in1(N__6308),
            .in2(_gnd_net_),
            .in3(N__8125),
            .lcout(\U712_CHIP_RAM.N_555 ),
            .ltout(\U712_CHIP_RAM.N_555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_11_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_11_7_5 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_2_LC_11_7_5  (
            .in0(N__7981),
            .in1(_gnd_net_),
            .in2(N__6182),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER16 ),
            .ltout(\U712_CHIP_RAM.SDRAM_COUNTER16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DBENn_LC_11_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBENn_LC_11_7_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBENn_LC_11_7_6 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \U712_CHIP_RAM.DBENn_LC_11_7_6  (
            .in0(N__6173),
            .in1(N__11046),
            .in2(N__6164),
            .in3(N__8432),
            .lcout(DBENn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10236),
            .ce(),
            .sr(N__10680));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_11_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_11_8_0 .LUT_INIT=16'b1101111111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIKHPV5_2_LC_11_8_0  (
            .in0(N__6457),
            .in1(N__8005),
            .in2(N__6380),
            .in3(N__10547),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERe_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_11_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_11_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_11_8_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNO_0_LC_11_8_1  (
            .in0(N__6364),
            .in1(N__7378),
            .in2(_gnd_net_),
            .in3(N__7683),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_11_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_11_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIOV791_LC_11_8_2  (
            .in0(N__7580),
            .in1(N__8004),
            .in2(_gnd_net_),
            .in3(N__8118),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_355_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_11_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_11_8_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIL6NI4_LC_11_8_3  (
            .in0(N__10546),
            .in1(N__7377),
            .in2(N__6341),
            .in3(N__7682),
            .lcout(\U712_CHIP_RAM.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_11_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_11_8_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_3_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__7873),
            .in2(_gnd_net_),
            .in3(N__7285),
            .lcout(\U712_CHIP_RAM.N_289 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_11_8_5  (
            .in0(N__8007),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6456),
            .lcout(\U712_CHIP_RAM.N_387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_3_LC_11_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_3_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_3_LC_11_8_6 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNITERT_0_3_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__7872),
            .in2(_gnd_net_),
            .in3(N__7286),
            .lcout(\U712_CHIP_RAM.N_293 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_11_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_11_8_7 .LUT_INIT=16'b0100010000001010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNILL5O1_0_LC_11_8_7  (
            .in0(N__8006),
            .in1(N__8119),
            .in2(N__7308),
            .in3(N__7581),
            .lcout(\U712_CHIP_RAM.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_11_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_11_9_0 .LUT_INIT=16'b0111011111110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNILE372_LC_11_9_0  (
            .in0(N__8116),
            .in1(N__8000),
            .in2(N__6317),
            .in3(N__7570),
            .lcout(\U712_CHIP_RAM.N_356 ),
            .ltout(\U712_CHIP_RAM.N_356_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_11_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_11_9_1 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_2_LC_11_9_1  (
            .in0(N__7875),
            .in1(N__7291),
            .in2(N__6512),
            .in3(N__7677),
            .lcout(\U712_CHIP_RAM.N_448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_9_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIAENR1_7_LC_11_9_2  (
            .in0(N__7801),
            .in1(N__7816),
            .in2(N__7754),
            .in3(N__7831),
            .lcout(\U712_CHIP_RAM.N_288 ),
            .ltout(\U712_CHIP_RAM.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_11_9_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_11_9_3 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNI3M1M2_LC_11_9_3  (
            .in0(N__7569),
            .in1(_gnd_net_),
            .in2(N__6503),
            .in3(N__8115),
            .lcout(\U712_CHIP_RAM.N_473 ),
            .ltout(\U712_CHIP_RAM.N_473_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_3_LC_11_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_3_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_3_LC_11_9_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI05TJ3_3_LC_11_9_4  (
            .in0(N__7290),
            .in1(_gnd_net_),
            .in2(N__6488),
            .in3(N__7874),
            .lcout(\U712_CHIP_RAM.N_557 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_9_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_9_5 .LUT_INIT=16'b0001001100010100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_11_9_5  (
            .in0(N__7876),
            .in1(N__7293),
            .in2(N__7592),
            .in3(N__8117),
            .lcout(\U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_57_i_a2_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_9_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_9_6 .LUT_INIT=16'b0111001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_WRITE_CYCLE_LC_11_9_6  (
            .in0(N__6422),
            .in1(N__7040),
            .in2(N__11670),
            .in3(N__10509),
            .lcout(DMA_WRITE_CYCLE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10241),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5F93_0_LC_11_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5F93_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5F93_0_LC_11_9_7 .LUT_INIT=16'b1111111101011101;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIS5F93_0_LC_11_9_7  (
            .in0(N__10510),
            .in1(N__7292),
            .in2(N__8034),
            .in3(N__7678),
            .lcout(\U712_CHIP_RAM.N_362 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_LC_11_10_0  (
            .in0(N__6996),
            .in1(N__8040),
            .in2(_gnd_net_),
            .in3(N__6461),
            .lcout(DMA_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10249),
            .ce(N__6431),
            .sr(N__10668));
    defparam \U712_CHIP_RAM.DBDIR_LC_11_11_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_11_6 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.DBDIR_LC_11_11_6 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \U712_CHIP_RAM.DBDIR_LC_11_11_6  (
            .in0(N__7032),
            .in1(N__6391),
            .in2(_gnd_net_),
            .in3(N__6421),
            .lcout(DBDIR_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10252),
            .ce(),
            .sr(N__10666));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_LC_11_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_LC_11_12_1 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_LC_11_12_1  (
            .in0(N__11163),
            .in1(N__11748),
            .in2(_gnd_net_),
            .in3(N__11062),
            .lcout(\U712_BYTE_ENABLE.N_451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_7 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \U712_CHIP_RAM.CAS_SYNC_0_LC_11_12_7  (
            .in0(N__10486),
            .in1(N__9901),
            .in2(_gnd_net_),
            .in3(N__11749),
            .lcout(\U712_CHIP_RAM.CAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10256),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_13_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_13_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_1_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__9370),
            .in2(_gnd_net_),
            .in3(N__8294),
            .lcout(),
            .ltout(\U712_REG_SM.N_306_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_13_1 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_1_LC_11_13_1 .LUT_INIT=16'b1110000000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_1_LC_11_13_1  (
            .in0(N__8337),
            .in1(N__6619),
            .in2(N__6599),
            .in3(N__10491),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10259),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_4 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_4 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \U712_REG_SM.REG_CYCLE_RNO_0_LC_11_13_4  (
            .in0(N__8228),
            .in1(N__6586),
            .in2(N__9380),
            .in3(N__6573),
            .lcout(),
            .ltout(\U712_REG_SM.N_399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_CYCLE_LC_11_13_5 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_REG_SM.REG_CYCLE_LC_11_13_5  (
            .in0(N__10113),
            .in1(N__10490),
            .in2(N__6596),
            .in3(N__6593),
            .lcout(REG_CYCLEm),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10259),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_6 .LUT_INIT=16'b1010100011111101;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNO_0_2_LC_11_13_6  (
            .in0(N__8336),
            .in1(N__8295),
            .in2(N__9379),
            .in3(N__6574),
            .lcout(),
            .ltout(\U712_REG_SM.N_353_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_2_LC_11_13_7 .LUT_INIT=16'b0000101100000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_2_LC_11_13_7  (
            .in0(N__6587),
            .in1(N__9377),
            .in2(N__6578),
            .in3(N__10492),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10259),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.C3_SYNC_1_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.C3_SYNC_1_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6557),
            .lcout(\U712_REG_SM.C3_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10263),
            .ce(),
            .sr(N__10662));
    defparam \U712_REG_SM.REG_TACK_LC_11_14_2 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.REG_TACK_LC_11_14_2 .LUT_INIT=16'b1111111000010000;
    LogicCell40 \U712_REG_SM.REG_TACK_LC_11_14_2  (
            .in0(N__6680),
            .in1(N__6707),
            .in2(N__6540),
            .in3(N__6548),
            .lcout(REG_TACK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10263),
            .ce(),
            .sr(N__10662));
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_14_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_14_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.STATE_COUNT_0_LC_11_14_7 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_0_LC_11_14_7  (
            .in0(N__6743),
            .in1(N__6695),
            .in2(_gnd_net_),
            .in3(N__8225),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10263),
            .ce(),
            .sr(N__10662));
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_1 .C_ON=1'b0;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_1 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \U712_REG_SM.REG_TACK_RNO_1_LC_11_15_1  (
            .in0(N__6730),
            .in1(N__6661),
            .in2(N__8226),
            .in3(N__6693),
            .lcout(\U712_REG_SM.un1_STATE_COUNT_3_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_2 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_5_LC_11_15_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_5_LC_11_15_2  (
            .in0(N__10505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6668),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.LDSn_RNO_0_LC_11_15_3 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \U712_REG_SM.LDSn_RNO_0_LC_11_15_3  (
            .in0(N__11534),
            .in1(N__11375),
            .in2(N__9809),
            .in3(N__11465),
            .lcout(\U712_REG_SM.N_432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_15_4 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_7_LC_11_15_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_7_LC_11_15_4  (
            .in0(N__10507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6653),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_15_5 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_8_LC_11_15_5 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_8_LC_11_15_5  (
            .in0(N__6701),
            .in1(N__10508),
            .in2(N__8227),
            .in3(N__6694),
            .lcout(\U712_REG_SM.STATE_COUNTZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_6 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_6 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_4_LC_11_15_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_4_LC_11_15_6  (
            .in0(N__10504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6679),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_15_7 .SEQ_MODE=4'b1000;
    defparam \U712_REG_SM.STATE_COUNT_6_LC_11_15_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_REG_SM.STATE_COUNT_6_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(N__10506),
            .in2(_gnd_net_),
            .in3(N__6662),
            .lcout(\U712_REG_SM.STATE_COUNTZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10266),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_130_i_LC_11_19_5 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_130_i_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_130_i_LC_11_19_5 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \U712_BUFFERS.N_130_i_LC_11_19_5  (
            .in0(N__11677),
            .in1(N__9894),
            .in2(_gnd_net_),
            .in3(N__11750),
            .lcout(N_130_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_1_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_1_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WEn_LC_12_4_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WEn_LC_12_4_7 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.WEn_LC_12_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.WEn_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6902),
            .lcout(WEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10226),
            .ce(),
            .sr(N__10694));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_0 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_12_5_0  (
            .in0(N__10010),
            .in1(N__9217),
            .in2(N__6839),
            .in3(N__8810),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_12_5_2  (
            .in0(N__6830),
            .in1(N__6776),
            .in2(_gnd_net_),
            .in3(N__9216),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3 .LUT_INIT=16'b1111000111100000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_12_5_3  (
            .in0(N__9218),
            .in1(N__10012),
            .in2(N__6818),
            .in3(N__8801),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_12_5_5  (
            .in0(N__9215),
            .in1(N__6815),
            .in2(_gnd_net_),
            .in3(N__7124),
            .lcout(),
            .ltout(\U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6 .LUT_INIT=16'b1111000011100100;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_12_5_6  (
            .in0(N__10011),
            .in1(N__8780),
            .in2(N__6800),
            .in3(N__9219),
            .lcout(\U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_12_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_12_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_12_5_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_4_LC_12_5_7  (
            .in0(N__6797),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10227),
            .ce(N__7060),
            .sr(N__10686));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_12_6_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_12_6_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_12_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_0_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6770),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_12_6_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_12_6_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_12_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_1_LC_12_6_1  (
            .in0(N__7238),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_12_6_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_12_6_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_12_6_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_2_LC_12_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7202),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_12_6_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_12_6_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_12_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_5_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7175),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_12_6_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_12_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_6_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7145),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_12_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_12_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_12_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_7_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7118),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_12_6_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_12_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \U712_CHIP_RAM.CPU_COL_ADDRESS_esr_3_LC_12_6_7  (
            .in0(N__7085),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\U712_CHIP_RAM.CPU_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10228),
            .ce(N__7064),
            .sr(N__10679));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_12_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_12_7_0 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_LC_12_7_0  (
            .in0(N__7036),
            .in1(N__9821),
            .in2(_gnd_net_),
            .in3(N__6998),
            .lcout(\U712_CHIP_RAM.WRITE_CYCLEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10231),
            .ce(N__6929),
            .sr(N__10673));
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI324S_LC_12_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI324S_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.DMA_CYCLE_esr_RNI324S_LC_12_8_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_CYCLE_esr_RNI324S_LC_12_8_0  (
            .in0(N__7983),
            .in1(N__11153),
            .in2(_gnd_net_),
            .in3(N__7600),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_294_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_12_8_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_12_8_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNI8MK44_1_LC_12_8_1  (
            .in0(N__8114),
            .in1(N__7374),
            .in2(N__7706),
            .in3(N__7686),
            .lcout(),
            .ltout(\U712_CHIP_RAM.N_469_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVM119_1_LC_12_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVM119_1_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNIVM119_1_LC_12_8_2 .LUT_INIT=16'b1111101111110011;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNIVM119_1_LC_12_8_2  (
            .in0(N__7419),
            .in1(N__10428),
            .in2(N__7631),
            .in3(N__7622),
            .lcout(\U712_CHIP_RAM.N_309 ),
            .ltout(\U712_CHIP_RAM.N_309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIUJS3D_LC_12_8_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIUJS3D_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIUJS3D_LC_12_8_3 .LUT_INIT=16'b1111100011111100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIUJS3D_LC_12_8_3  (
            .in0(N__7601),
            .in1(N__7514),
            .in2(N__7508),
            .in3(N__7984),
            .lcout(\U712_CHIP_RAM.N_200 ),
            .ltout(\U712_CHIP_RAM.N_200_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_8_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_8_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_8_4 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_12_8_4  (
            .in0(N__7247),
            .in1(N__7505),
            .in2(N__7499),
            .in3(N__7496),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10235),
            .ce(N__7739),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_8_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_8_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_8_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_12_8_5  (
            .in0(N__10427),
            .in1(N__7490),
            .in2(N__7919),
            .in3(N__7783),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10235),
            .ce(N__7739),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_12_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_12_8_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \U712_CHIP_RAM.WRITE_CYCLE_esr_RNI1IJO_LC_12_8_6  (
            .in0(N__7982),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7442),
            .lcout(\U712_CHIP_RAM.N_285 ),
            .ltout(\U712_CHIP_RAM.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_3_LC_12_8_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_3_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.CLK_EN_ess_RNO_3_LC_12_8_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \U712_CHIP_RAM.CLK_EN_ess_RNO_3_LC_12_8_7  (
            .in0(N__8113),
            .in1(N__10016),
            .in2(N__7388),
            .in3(N__7375),
            .lcout(\U712_CHIP_RAM.un1_SDRAM_COUNTER47_2_0_a2_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_12_9_0 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_12_9_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__7307),
            .in2(_gnd_net_),
            .in3(N__7241),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_0 ),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_12_9_1 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_12_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_12_9_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_12_9_1  (
            .in0(N__7784),
            .in1(N__8120),
            .in2(_gnd_net_),
            .in3(N__8054),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_0 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_12_9_2 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_12_9_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__8016),
            .in2(_gnd_net_),
            .in3(N__7910),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTER_s_2 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_1 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_9_3 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_9_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_9_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_12_9_3  (
            .in0(N__7785),
            .in1(N__7888),
            .in2(_gnd_net_),
            .in3(N__7835),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_2 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_9_4 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_9_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_12_9_4  (
            .in0(N__7781),
            .in1(N__7832),
            .in2(_gnd_net_),
            .in3(N__7820),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_3 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_12_9_5 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_12_9_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_12_9_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_12_9_5  (
            .in0(N__7786),
            .in1(N__7817),
            .in2(_gnd_net_),
            .in3(N__7805),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_4 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_12_9_6 .C_ON=1'b1;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_12_9_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_12_9_6  (
            .in0(N__7782),
            .in1(N__7802),
            .in2(_gnd_net_),
            .in3(N__7790),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6 ),
            .ltout(),
            .carryin(\U712_CHIP_RAM.SDRAM_COUNTER_cry_5 ),
            .carryout(\U712_CHIP_RAM.SDRAM_COUNTER_cry_6 ),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_12_9_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_12_9_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_12_9_7  (
            .in0(N__7787),
            .in1(N__7753),
            .in2(_gnd_net_),
            .in3(N__7757),
            .lcout(\U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10237),
            .ce(N__7732),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_12_10_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_12_10_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_1_LC_12_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_1_LC_12_10_0  (
            .in0(N__10424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10286),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10239),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_10_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_3_LC_12_10_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_3_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__10426),
            .in2(_gnd_net_),
            .in3(N__8405),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10239),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_12_10_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_2_LC_12_10_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_2_LC_12_10_6  (
            .in0(N__10425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8411),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10239),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_211_i_LC_12_12_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_211_i_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_211_i_LC_12_12_5 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \U712_BYTE_ENABLE.N_211_i_LC_12_12_5  (
            .in0(N__8351),
            .in1(N__11610),
            .in2(N__9395),
            .in3(N__8399),
            .lcout(N_211_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_12_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_12_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_1_LC_12_12_6  (
            .in0(N__11744),
            .in1(N__11164),
            .in2(_gnd_net_),
            .in3(N__11078),
            .lcout(),
            .ltout(\U712_BYTE_ENABLE.N_410_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_148_i_LC_12_12_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_148_i_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_148_i_LC_12_12_7 .LUT_INIT=16'b0000000000001101;
    LogicCell40 \U712_BYTE_ENABLE.N_148_i_LC_12_12_7  (
            .in0(N__8350),
            .in1(N__11609),
            .in2(N__8372),
            .in3(N__9391),
            .lcout(N_148_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_12_13_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_12_13_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLLBEn_i_a2_0_0_LC_12_13_0  (
            .in0(N__10069),
            .in1(N__11530),
            .in2(_gnd_net_),
            .in3(N__11379),
            .lcout(\U712_BYTE_ENABLE.un1_CLLBEn_i_a2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_12_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_12_14_0 .LUT_INIT=16'b0000111000000010;
    LogicCell40 \U712_REG_SM.STATE_COUNT_RNI3HF31_1_LC_12_14_0  (
            .in0(N__8329),
            .in1(N__9345),
            .in2(N__8296),
            .in3(N__8213),
            .lcout(\U712_REG_SM.N_95 ),
            .ltout(\U712_REG_SM.N_95_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_1 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.ASn_ess_RNO_LC_12_14_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \U712_REG_SM.ASn_ess_RNO_LC_12_14_1  (
            .in0(N__10729),
            .in1(_gnd_net_),
            .in2(N__8183),
            .in3(_gnd_net_),
            .lcout(\U712_REG_SM.N_95_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.LDSn_LC_12_15_3 .C_ON=1'b0;
    defparam \U712_REG_SM.LDSn_LC_12_15_3 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.LDSn_LC_12_15_3 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \U712_REG_SM.LDSn_LC_12_15_3  (
            .in0(N__8164),
            .in1(N__8681),
            .in2(N__9378),
            .in3(N__8180),
            .lcout(LDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10261),
            .ce(),
            .sr(N__10657));
    defparam \U712_REG_SM.UDSn_LC_12_15_7 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_LC_12_15_7 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.UDSn_LC_12_15_7 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \U712_REG_SM.UDSn_LC_12_15_7  (
            .in0(N__8642),
            .in1(N__8680),
            .in2(N__8659),
            .in3(N__9369),
            .lcout(UDSn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10261),
            .ce(),
            .sr(N__10657));
    defparam \U712_REG_SM.UDSn_RNO_0_LC_12_16_1 .C_ON=1'b0;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \U712_REG_SM.UDSn_RNO_0_LC_12_16_1 .LUT_INIT=16'b0000010001000000;
    LogicCell40 \U712_REG_SM.UDSn_RNO_0_LC_12_16_1  (
            .in0(N__9810),
            .in1(N__11506),
            .in2(N__11381),
            .in3(N__11466),
            .lcout(\U712_REG_SM.N_433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_1.C_ON=1'b0;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_1.SEQ_MODE=4'b0000;
    defparam RESETn_ibuf_RNIM9SF_LC_12_19_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 RESETn_ibuf_RNIM9SF_LC_12_19_1 (
            .in0(N__10469),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(RESETn_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_5_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_5_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_3_LC_13_5_3 .LUT_INIT=16'b1100100001000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_3_LC_13_5_3  (
            .in0(N__8504),
            .in1(N__8580),
            .in2(N__8627),
            .in3(N__9563),
            .lcout(CMA_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10230),
            .ce(N__11218),
            .sr(N__10696));
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_4_LC_13_5_4 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_4_LC_13_5_4  (
            .in0(N__8581),
            .in1(N__8438),
            .in2(N__8520),
            .in3(N__8603),
            .lcout(CMA_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10230),
            .ce(N__11218),
            .sr(N__10696));
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_6_LC_13_5_7 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_6_LC_13_5_7  (
            .in0(N__8582),
            .in1(N__9677),
            .in2(N__8519),
            .in3(N__8465),
            .lcout(CMA_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10230),
            .ce(N__11218),
            .sr(N__10696));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_6_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_13_6_6  (
            .in0(N__9655),
            .in1(N__10996),
            .in2(_gnd_net_),
            .in3(N__9065),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10793),
            .ce(N__10766),
            .sr(N__10689));
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_7_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_7_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_A1_nesr_LC_13_7_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_A1_nesr_LC_13_7_0  (
            .in0(N__10982),
            .in1(N__8967),
            .in2(_gnd_net_),
            .in3(N__8927),
            .lcout(\U712_CHIP_RAM.DMA_AZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_7_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_7_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_7_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_7_1  (
            .in0(N__8968),
            .in1(N__10983),
            .in2(_gnd_net_),
            .in3(N__9022),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_2 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_7_2  (
            .in0(N__9023),
            .in1(_gnd_net_),
            .in2(N__10998),
            .in3(N__9599),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_7_4 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_13_7_4  (
            .in0(N__9062),
            .in1(_gnd_net_),
            .in2(N__10999),
            .in3(N__9656),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_7_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_7_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_7_5  (
            .in0(N__9708),
            .in1(N__10990),
            .in2(_gnd_net_),
            .in3(N__9063),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_7_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_7_6  (
            .in0(N__9748),
            .in1(_gnd_net_),
            .in2(N__11000),
            .in3(N__9709),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_7_7  (
            .in0(N__8873),
            .in1(N__10994),
            .in2(_gnd_net_),
            .in3(N__9749),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_A1_nesrC_net ),
            .ce(N__10764),
            .sr(N__10681));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_8_0  (
            .in0(N__9009),
            .in1(_gnd_net_),
            .in2(N__8969),
            .in3(N__10980),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10762),
            .sr(N__10674));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_13_8_6  (
            .in0(N__10846),
            .in1(N__10981),
            .in2(_gnd_net_),
            .in3(N__8872),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10790),
            .ce(N__10762),
            .sr(N__10674));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_0 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_13_9_0  (
            .in0(N__8853),
            .in1(N__10979),
            .in2(_gnd_net_),
            .in3(N__10845),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net ),
            .ce(N__10761),
            .sr(N__10672));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_7 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_8_LC_13_10_7  (
            .in0(N__8729),
            .in1(N__10945),
            .in2(N__10847),
            .in3(N__8698),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_8C_net ),
            .ce(),
            .sr(N__10669));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_13_13_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_13_13_6 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_a2_0_LC_13_13_6  (
            .in0(N__10070),
            .in1(N__11380),
            .in2(_gnd_net_),
            .in3(N__11470),
            .lcout(\U712_BYTE_ENABLE.N_409 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_REG_SM.ASn_ess_LC_13_14_0 .C_ON=1'b0;
    defparam \U712_REG_SM.ASn_ess_LC_13_14_0 .SEQ_MODE=4'b1001;
    defparam \U712_REG_SM.ASn_ess_LC_13_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_REG_SM.ASn_ess_LC_13_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9363),
            .lcout(ASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10264),
            .ce(N__9251),
            .sr(N__10663));
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_13_20_6 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.LLBE_0_LC_13_20_6 .LUT_INIT=16'b0000011101010000;
    LogicCell40 \U712_BYTE_ENABLE.LLBE_0_LC_13_20_6  (
            .in0(N__11611),
            .in1(N__11547),
            .in2(N__11362),
            .in3(N__11440),
            .lcout(LLBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CASn_LC_14_5_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_5 .SEQ_MODE=4'b1001;
    defparam \U712_CHIP_RAM.CASn_LC_14_5_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \U712_CHIP_RAM.CASn_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9227),
            .lcout(CASn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10234),
            .ce(),
            .sr(N__10702));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_6_5 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_6_5 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_6_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_6_5  (
            .in0(N__10995),
            .in1(N__9710),
            .in2(_gnd_net_),
            .in3(N__9064),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10792),
            .ce(N__10768),
            .sr(N__10697));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_14_7_2  (
            .in0(N__9016),
            .in1(N__10936),
            .in2(_gnd_net_),
            .in3(N__9595),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(N__10767),
            .sr(N__10690));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_3 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_3 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_14_7_3  (
            .in0(N__8955),
            .in1(N__10935),
            .in2(_gnd_net_),
            .in3(N__8926),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(N__10767),
            .sr(N__10690));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_7_4  (
            .in0(N__9747),
            .in1(N__10938),
            .in2(_gnd_net_),
            .in3(N__8871),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(N__10767),
            .sr(N__10690));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_7_6  (
            .in0(N__9746),
            .in1(N__10937),
            .in2(_gnd_net_),
            .in3(N__9699),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10791),
            .ce(N__10767),
            .sr(N__10690));
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_14_8_6  (
            .in0(N__10934),
            .in1(N__9651),
            .in2(_gnd_net_),
            .in3(N__9594),
            .lcout(\U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net ),
            .ce(N__10765),
            .sr(N__10682));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_9_4 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_9_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_9_4  (
            .in0(N__10933),
            .in1(N__9650),
            .in2(_gnd_net_),
            .in3(N__9593),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10789),
            .ce(N__10763),
            .sr(N__10675));
    defparam \U712_BYTE_ENABLE.N_146_i_LC_14_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_146_i_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_146_i_LC_14_12_1 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \U712_BYTE_ENABLE.N_146_i_LC_14_12_1  (
            .in0(N__9428),
            .in1(N__11089),
            .in2(N__9875),
            .in3(N__11172),
            .lcout(N_146_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam pll_RNI8MQ3_LC_14_12_5.C_ON=1'b0;
    defparam pll_RNI8MQ3_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam pll_RNI8MQ3_LC_14_12_5.LUT_INIT=16'b0101010101010101;
    LogicCell40 pll_RNI8MQ3_LC_14_12_5 (
            .in0(N__9529),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CLK40_PLL_i_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_0 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_0 .LUT_INIT=16'b0011000001110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUUBEn_i_a2_LC_14_13_0  (
            .in0(N__11621),
            .in1(N__9422),
            .in2(N__10090),
            .in3(N__11549),
            .lcout(\U712_BYTE_ENABLE.N_406 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_13_4 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_13_4 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \U712_BYTE_ENABLE.un1_CLMBEn_i_a2_LC_14_13_4  (
            .in0(N__11620),
            .in1(N__9421),
            .in2(N__10089),
            .in3(N__11548),
            .lcout(\U712_BYTE_ENABLE.N_411 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_14_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_14_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \U712_BYTE_ENABLE.un1_CUMBEn_i_x2_LC_14_14_1  (
            .in0(N__11471),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11336),
            .lcout(\U712_BYTE_ENABLE.N_284_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_374_i_LC_14_20_3 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_374_i_LC_14_20_3 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_374_i_LC_14_20_3 .LUT_INIT=16'b0000110111010000;
    LogicCell40 \U712_BYTE_ENABLE.N_374_i_LC_14_20_3  (
            .in0(N__11613),
            .in1(N__11551),
            .in2(N__11463),
            .in3(N__11349),
            .lcout(N_374_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.N_373_i_LC_14_20_5 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_373_i_LC_14_20_5 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_373_i_LC_14_20_5 .LUT_INIT=16'b0000111011100000;
    LogicCell40 \U712_BYTE_ENABLE.N_373_i_LC_14_20_5  (
            .in0(N__11612),
            .in1(N__11550),
            .in2(N__11462),
            .in3(N__11348),
            .lcout(N_373_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_7 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.UMBE_0_LC_14_20_7 .LUT_INIT=16'b0000101010110000;
    LogicCell40 \U712_BYTE_ENABLE.UMBE_0_LC_14_20_7  (
            .in0(N__11614),
            .in1(N__11552),
            .in2(N__11464),
            .in3(N__11350),
            .lcout(UMBEn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_7_6 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_7_6 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.CMA_esr_9_LC_15_7_6 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \U712_CHIP_RAM.CMA_esr_9_LC_15_7_6  (
            .in0(N__11270),
            .in1(N__11261),
            .in2(N__10079),
            .in3(N__10799),
            .lcout(CMA_c_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10242),
            .ce(N__11222),
            .sr(N__10698));
    defparam \U712_BYTE_ENABLE.N_150_i_LC_15_12_1 .C_ON=1'b0;
    defparam \U712_BYTE_ENABLE.N_150_i_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \U712_BYTE_ENABLE.N_150_i_LC_15_12_1 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \U712_BYTE_ENABLE.N_150_i_LC_15_12_1  (
            .in0(N__11173),
            .in1(N__11099),
            .in2(N__9902),
            .in3(N__11088),
            .lcout(N_150_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_2 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_2 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_16_8_2  (
            .in0(N__10309),
            .in1(N__10978),
            .in2(_gnd_net_),
            .in3(N__10832),
            .lcout(\U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10788),
            .ce(N__10769),
            .sr(N__10699));
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_1 .C_ON=1'b0;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \U712_CHIP_RAM.RAS_SYNC_0_LC_17_9_1  (
            .in0(N__10470),
            .in1(N__10325),
            .in2(_gnd_net_),
            .in3(N__10313),
            .lcout(\U712_CHIP_RAM.RAS_SYNCZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__10260),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.N_136_i_LC_24_19_1 .C_ON=1'b0;
    defparam \U712_BUFFERS.N_136_i_LC_24_19_1 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.N_136_i_LC_24_19_1 .LUT_INIT=16'b0011001000110000;
    LogicCell40 \U712_BUFFERS.N_136_i_LC_24_19_1  (
            .in0(N__9858),
            .in1(N__10133),
            .in2(N__10094),
            .in3(N__11731),
            .lcout(N_136_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3 .C_ON=1'b0;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3 .SEQ_MODE=4'b0000;
    defparam \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3 .LUT_INIT=16'b0010000001111111;
    LogicCell40 \U712_BUFFERS.DRDDIR_i_m2_LC_24_19_3  (
            .in0(N__9857),
            .in1(N__9820),
            .in2(N__11743),
            .in3(N__11687),
            .lcout(N_357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // U712_TOP

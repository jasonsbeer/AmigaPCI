-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jul 1 2025 18:43:57

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U409_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U409_TOP
entity U409_TOP is
port (
    ROM_DELAY : in std_logic_vector(1 downto 0);
    F_BANK : out std_logic_vector(1 downto 0);
    PCIAT : out std_logic_vector(1 downto 0);
    TM : in std_logic_vector(2 downto 0);
    TT : in std_logic_vector(1 downto 0);
    A : in std_logic_vector(31 downto 1);
    D : inout std_logic_vector(7 downto 4);
    PCS0 : out std_logic;
    F_ENn : out std_logic;
    TSn : in std_logic;
    SPIO_J : in std_logic;
    SPIO : out std_logic;
    RTC_ENn : out std_logic;
    RESETn : in std_logic;
    OVL : in std_logic;
    F_RDY : in std_logic;
    CONFIGENn : out std_logic;
    PPIO : out std_logic;
    PORTSIZE : out std_logic;
    F_RSTn : out std_logic;
    TICK60 : out std_logic;
    PCS1 : out std_logic;
    CIACS0n : out std_logic;
    SCS0 : out std_logic;
    CPUCONFn : in std_logic;
    CLK6 : in std_logic;
    AGNUS_CLK : out std_logic;
    CLK_CIA : out std_logic;
    BUFENn : out std_logic;
    AUTOBOOT : in std_logic;
    RnW : in std_logic;
    XCLK : in std_logic;
    F_WRITEn : out std_logic;
    F_READn : out std_logic;
    CIACS1n : out std_logic;
    PPIO_J : in std_logic;
    TICK50 : out std_logic;
    TCIn : out std_logic;
    TBIn : out std_logic;
    RAMSPACEn : out std_logic;
    BPRO_ENn : out std_logic;
    CLK40_IN : in std_logic;
    CLK28_IN : in std_logic;
    XCLK_ENn : in std_logic;
    SCS1 : out std_logic;
    REGSPACEn : out std_logic;
    F_WPn : out std_logic;
    ATA_ENn : out std_logic;
    TACKn : inout std_logic;
    BREG_ENn : out std_logic;
    ROMENn : out std_logic);
end U409_TOP;

-- Architecture of U409_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U409_TOP is

signal \N__13653\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13613\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13595\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13549\ : std_logic;
signal \N__13548\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13539\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13530\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13514\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13512\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13458\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13441\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13406\ : std_logic;
signal \N__13405\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13395\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13379\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13369\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13332\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13314\ : std_logic;
signal \N__13307\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13296\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13271\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13260\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13244\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13242\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13162\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13144\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13108\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13081\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13064\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13055\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13046\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13036\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13009\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13001\ : std_logic;
signal \N__13000\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12991\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12974\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12965\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12956\ : std_logic;
signal \N__12955\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12947\ : std_logic;
signal \N__12946\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12938\ : std_logic;
signal \N__12937\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12928\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12919\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12911\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12893\ : std_logic;
signal \N__12892\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12874\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12868\ : std_logic;
signal \N__12865\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12859\ : std_logic;
signal \N__12856\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12850\ : std_logic;
signal \N__12847\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12823\ : std_logic;
signal \N__12820\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12814\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12796\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12787\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12775\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12769\ : std_logic;
signal \N__12766\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12760\ : std_logic;
signal \N__12757\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12742\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12725\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12704\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12701\ : std_logic;
signal \N__12698\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12625\ : std_logic;
signal \N__12622\ : std_logic;
signal \N__12619\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12601\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12568\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12541\ : std_logic;
signal \N__12538\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12528\ : std_logic;
signal \N__12525\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12487\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12466\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12460\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12373\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12361\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12242\ : std_logic;
signal \N__12239\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12233\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12136\ : std_logic;
signal \N__12133\ : std_logic;
signal \N__12130\ : std_logic;
signal \N__12127\ : std_logic;
signal \N__12124\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11842\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11836\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11287\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11269\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10914\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10908\ : std_logic;
signal \N__10905\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10887\ : std_logic;
signal \N__10884\ : std_logic;
signal \N__10881\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10774\ : std_logic;
signal \N__10759\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10756\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10726\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10720\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10682\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10519\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10506\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10426\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10414\ : std_logic;
signal \N__10411\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10249\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10218\ : std_logic;
signal \N__10215\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10116\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10110\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9943\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9914\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9741\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9699\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9519\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9483\ : std_logic;
signal \N__9480\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9408\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9288\ : std_logic;
signal \N__9285\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9216\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9089\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8939\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8933\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8903\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8891\ : std_logic;
signal \N__8888\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8853\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8454\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8439\ : std_logic;
signal \N__8436\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8270\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8264\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8244\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8224\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8199\ : std_logic;
signal \N__8196\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8055\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8040\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8030\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8000\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7989\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7983\ : std_logic;
signal \N__7980\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7943\ : std_logic;
signal \N__7940\ : std_logic;
signal \N__7937\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7906\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7890\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7881\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7866\ : std_logic;
signal \N__7865\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7847\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7809\ : std_logic;
signal \N__7806\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7746\ : std_logic;
signal \N__7743\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7724\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7710\ : std_logic;
signal \N__7707\ : std_logic;
signal \N__7704\ : std_logic;
signal \N__7701\ : std_logic;
signal \N__7698\ : std_logic;
signal \N__7695\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7686\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7670\ : std_logic;
signal \N__7667\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7653\ : std_logic;
signal \N__7650\ : std_logic;
signal \N__7647\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7635\ : std_logic;
signal \N__7632\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7626\ : std_logic;
signal \N__7625\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7614\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7608\ : std_logic;
signal \N__7605\ : std_logic;
signal \N__7602\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7560\ : std_logic;
signal \N__7557\ : std_logic;
signal \N__7554\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7542\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7530\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7512\ : std_logic;
signal \N__7509\ : std_logic;
signal \N__7506\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7485\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7471\ : std_logic;
signal \N__7468\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7452\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7449\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7437\ : std_logic;
signal \N__7436\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7397\ : std_logic;
signal \N__7394\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7359\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7338\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7284\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7260\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7252\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7242\ : std_logic;
signal \N__7233\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7227\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7224\ : std_logic;
signal \N__7221\ : std_logic;
signal \N__7218\ : std_logic;
signal \N__7215\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7191\ : std_logic;
signal \N__7188\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7172\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7155\ : std_logic;
signal \N__7152\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7116\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7107\ : std_logic;
signal \N__7104\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7074\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7017\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6954\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6945\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6912\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6894\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6882\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6876\ : std_logic;
signal \N__6873\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6864\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6849\ : std_logic;
signal \N__6846\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6813\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6776\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6702\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6666\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6539\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6480\ : std_logic;
signal \N__6477\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6429\ : std_logic;
signal \N__6426\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6381\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6375\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6348\ : std_logic;
signal \N__6345\ : std_logic;
signal \N__6342\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6264\ : std_logic;
signal \N__6261\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6246\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6237\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5985\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5919\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5862\ : std_logic;
signal \N__5859\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5727\ : std_logic;
signal \N__5724\ : std_logic;
signal \N__5721\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5715\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5691\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5670\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5661\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5613\ : std_logic;
signal \N__5610\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5514\ : std_logic;
signal \N__5511\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5505\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5493\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5304\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5271\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5163\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5103\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5097\ : std_logic;
signal \N__5094\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5052\ : std_logic;
signal \N__5049\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4995\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4947\ : std_logic;
signal \N__4944\ : std_logic;
signal \N__4941\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4867\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4854\ : std_logic;
signal \N__4851\ : std_logic;
signal \N__4846\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4818\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4812\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4723\ : std_logic;
signal \CLK80_OUT\ : std_logic;
signal \PPIO_c\ : std_logic;
signal \GNDG0\ : std_logic;
signal \SPIO_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \A_c_27\ : std_logic;
signal \A_c_28\ : std_logic;
signal \A_c_26\ : std_logic;
signal \U409_ADDRESS_DECODE.m12Z0Z_5\ : std_logic;
signal \U409_ADDRESS_DECODE.m12Z0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_13Z0Z_1\ : std_logic;
signal \A_c_25\ : std_logic;
signal \A_c_24\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_BPRO_ENn_i\ : std_logic;
signal \A_c_29\ : std_logic;
signal \U409_ADDRESS_DECODE.N_26_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.m54Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.un1_A_13Z0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0\ : std_logic;
signal \A_c_30\ : std_logic;
signal \A_c_31\ : std_logic;
signal \U409_ADDRESS_DECODE.N_59\ : std_logic;
signal \U409_ADDRESS_DECODE.N_59_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\ : std_logic;
signal \TT_c_1\ : std_logic;
signal \TT_c_0\ : std_logic;
signal \TM_c_2\ : std_logic;
signal \D_1_i\ : std_logic;
signal \CONFIGENn_c\ : std_logic;
signal \INVU409_AUTOCONFIG.CONFIGENnC_net\ : std_logic;
signal \PRO_BASE_2\ : std_logic;
signal \PRO_BASE_0\ : std_logic;
signal \PRO_BASE_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_CONFC_net\ : std_logic;
signal \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0\ : std_logic;
signal \U409_AUTOCONFIG.N_216_3_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_108\ : std_logic;
signal \U409_AUTOCONFIG.N_108_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_8\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_9\ : std_logic;
signal \U409_ADDRESS_DECODE_AUTOVECTOR_10\ : std_logic;
signal \U409_AUTOCONFIG.N_99\ : std_logic;
signal \U409_AUTOCONFIG.N_100\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\ : std_logic;
signal \D_OUT_2\ : std_logic;
signal \D_OUT_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_111\ : std_logic;
signal \U409_AUTOCONFIG.N_105_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_91\ : std_logic;
signal \U409_AUTOCONFIG.N_91_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\ : std_logic;
signal \INVU409_AUTOCONFIG.PR_OUT_1C_net\ : std_logic;
signal \U409_AUTOCONFIG.N_216_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.N_116\ : std_logic;
signal \U409_AUTOCONFIG.N_89\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_2\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\ : std_logic;
signal \PORTSIZE_0_i\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_6\ : std_logic;
signal \U409_AUTOCONFIG.N_109_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_117\ : std_logic;
signal \U409_AUTOCONFIG.N_113\ : std_logic;
signal \AUTOBOOT_c\ : std_logic;
signal \U409_AUTOCONFIG.N_101\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_119\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.D_OUT_sm0_0_cascade_\ : std_logic;
signal \D_OUT_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.PR_OUTZ0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.D_OUT_sm0_0\ : std_logic;
signal \D_OUT_0\ : std_logic;
signal \U409_AUTOCONFIG.N_90\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.N_98\ : std_logic;
signal \CPUCONFn_c\ : std_logic;
signal \U409_AUTOCONFIG.STATE4_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.N_104\ : std_logic;
signal \U409_AUTOCONFIG.N_103_cascade_\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\ : std_logic;
signal \A_c_4\ : std_logic;
signal \A_c_2\ : std_logic;
signal \U409_AUTOCONFIG.N_109\ : std_logic;
signal \U409_AUTOCONFIG.N_115\ : std_logic;
signal \U409_AUTOCONFIG.AC_STARTZ0\ : std_logic;
signal \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\ : std_logic;
signal \U409_CIA.CLK_CIA_r_1_0_cascade_\ : std_logic;
signal \bfn_8_12_0_\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_1\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_2\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_3\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_4\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_5\ : std_logic;
signal \U409_CIA.un2_CIA_CLK_COUNT_cry_6\ : std_logic;
signal \U409_CIA.CLK_CIA6_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn_i\ : std_logic;
signal \BRIDGE_BASE_2\ : std_logic;
signal \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\ : std_logic;
signal \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net\ : std_logic;
signal \BRIDGE_BASE_0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_BREG_ENn_i\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONFZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0\ : std_logic;
signal \BRIDGE_BASE_4\ : std_logic;
signal \BRIDGE_BASE_7\ : std_logic;
signal \A_c_7\ : std_logic;
signal \A_c_5\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6Z0Z_1\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6_0\ : std_logic;
signal \A_c_1\ : std_logic;
signal \U409_AUTOCONFIG.un1_STATE_6_0_cascade_\ : std_logic;
signal \D_in_6\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_\ : std_logic;
signal \BRIDGE_BASE_6\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\ : std_logic;
signal \CIA_SPACE\ : std_logic;
signal \U409_CIA.VMA_RNOZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn_i\ : std_logic;
signal \U409_CIA.un1_CIA_CLK_COUNT_3_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_2\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_5\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_3\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_4\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11_3_cascade_\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNT11\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_0\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_1\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_7\ : std_logic;
signal \U409_CIA.CIA_CLK_COUNTZ0Z_6\ : std_logic;
signal \U409_CIA.CLK_CIA6_4\ : std_logic;
signal \U409_ADDRESS_DECODE.N_77_mux_cascade_\ : std_logic;
signal \N_22_0_i\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RTC_ENn\ : std_logic;
signal \U409_ADDRESS_DECODE.PORTSIZE_2\ : std_logic;
signal \A_c_18\ : std_logic;
signal \LIDE_BASE_1\ : std_logic;
signal \A_c_17\ : std_logic;
signal \LIDE_BASE_2\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\ : std_logic;
signal \CONFIGURED\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\ : std_logic;
signal \LIDE_BASE_6\ : std_logic;
signal \LIDE_BASE_5\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0\ : std_logic;
signal \BRIDGE_BASE_5\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0\ : std_logic;
signal \U409_AUTOCONFIG.un1_AZ0Z_13\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONFZ0\ : std_logic;
signal \D_in_5\ : std_logic;
signal \BRIDGE_BASE_1\ : std_logic;
signal \LIDE_BASE_7\ : std_logic;
signal \D_in_7\ : std_logic;
signal \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1\ : std_logic;
signal \BRIDGE_BASE_3\ : std_logic;
signal \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1\ : std_logic;
signal \D_in_4\ : std_logic;
signal \un1_AUTOCONFIG_SPACE\ : std_logic;
signal \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\ : std_logic;
signal \N_71_mux_cascade_\ : std_logic;
signal \N_23_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.m33Z0Z_3\ : std_logic;
signal \U409_ADDRESS_DECODE.m27Z0Z_3_cascade_\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4\ : std_logic;
signal \U409_ADDRESS_DECODE_m33_1\ : std_logic;
signal \U409_ADDRESS_DECODE_m33_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\ : std_logic;
signal \N_23\ : std_logic;
signal \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_4\ : std_logic;
signal \U409_ADDRESS_DECODE.CIA_SPACE_5\ : std_logic;
signal \LIDE_BASE_4\ : std_logic;
signal \LIDE_BASE_3\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\ : std_logic;
signal \AUTOCONFIG_SPACE\ : std_logic;
signal \BUFENn_c\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_SPACEZ0\ : std_logic;
signal \U409_ADDRESS_DECODE.ATA_ENZ0\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_ATA_ENn_i\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7\ : std_logic;
signal \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\ : std_logic;
signal \U409_AUTOCONFIG.STATE4\ : std_logic;
signal \INVU409_AUTOCONFIG.STATE_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\ : std_logic;
signal \N_71_mux\ : std_logic;
signal \N_70_mux\ : std_logic;
signal \U409_TRANSFER_ACK.N_20_0\ : std_logic;
signal \U409_AUTOCONFIG.STATE_d_2\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_1\ : std_logic;
signal \RnW_c\ : std_logic;
signal \U409_AUTOCONFIG.STATEZ0Z_0\ : std_logic;
signal \INVU409_AUTOCONFIG.AC_TACKC_net\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_REGSPACEn\ : std_logic;
signal \TACKn_in\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\ : std_logic;
signal \GB_BUFFER_CLK40_IN_c_g_THRU_CO\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_13\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS1n_i\ : std_logic;
signal \CIA_ENABLE\ : std_logic;
signal \CIA_ENABLE_cascade_\ : std_logic;
signal \A_c_12\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_CIACS0n_i\ : std_logic;
signal \U409_ADDRESS_DECODE.N_75\ : std_logic;
signal \N_77_mux_i\ : std_logic;
signal \U409_ADDRESS_DECODE.N_60_1\ : std_logic;
signal \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\ : std_logic;
signal \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\ : std_logic;
signal \AC_TACK\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.TACK_COUNTER6\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\ : std_logic;
signal \U409_ADDRESS_DECODE.Z2_SPACE\ : std_logic;
signal \ROMEN_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_\ : std_logic;
signal \U409_ADDRESS_DECODE.un1_RTC_ENn_2\ : std_logic;
signal \U409_ADDRESS_DECODE.N_61\ : std_logic;
signal \U409_TRANSFER_ACK.N_42_i_cascade_\ : std_logic;
signal \A_c_23\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1\ : std_logic;
signal \A_c_19\ : std_logic;
signal \A_c_22\ : std_logic;
signal \OVL_c\ : std_logic;
signal \A_c_21\ : std_logic;
signal \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\ : std_logic;
signal \ROMEN\ : std_logic;
signal \TACK_EN\ : std_logic;
signal \TCIn_1_i\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_ENZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0\ : std_logic;
signal \ROMENn_c\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROMENnC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_42_i\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\ : std_logic;
signal \PCIAT_c_1\ : std_logic;
signal \TM_c_0\ : std_logic;
signal \U409_ADDRESS_DECODE.N_58_mux\ : std_logic;
signal \TM_c_1\ : std_logic;
signal \PCIAT_c_0\ : std_logic;
signal \bfn_14_6_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_1\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_2\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_3\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_4\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_5\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_6\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_7\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_8\ : std_logic;
signal \bfn_14_7_0_\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_9\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_10\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_11\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_12\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_13\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_14\ : std_logic;
signal \U409_TICK.un3_COUNTER60_1_cry_15\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_TACK_ENZ0\ : std_logic;
signal \U409_CIA.VMAZ0\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\ : std_logic;
signal \U409_TRANSFER_ACK.N_33\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0\ : std_logic;
signal \ROM_DELAY_c_0\ : std_logic;
signal \ROM_DELAY_c_1\ : std_logic;
signal \U409_TRANSFER_ACK.N_31_i\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_4\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_8\ : std_logic;
signal \U409_TICK.TICK603_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_10\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_7\ : std_logic;
signal \U409_TICK.TICK603_10_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_0\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_12\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_2\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_16\ : std_logic;
signal \U409_TICK.TICK603_8\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_11\ : std_logic;
signal \U409_TICK.TICK603_11_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_3\ : std_logic;
signal \U409_TICK.TICK603_14_cascade_\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER60_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER60Z0Z_15\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\ : std_logic;
signal \CLK40_IN_c_g\ : std_logic;
signal \U409_TRANSFER_ACK.N_17_mux\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_3_0\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\ : std_logic;
signal \U409_TRANSFER_ACK.N_55_cascade_\ : std_logic;
signal \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\ : std_logic;
signal \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_1\ : std_logic;
signal \CLK_CIA_c\ : std_logic;
signal \U409_TRANSFER_ACK.LASTCLKZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.LASTCLK_1C_net\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0\ : std_logic;
signal \N_52_1\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\ : std_logic;
signal \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\ : std_logic;
signal \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \U409_TICK.TICK503_10_cascade_\ : std_logic;
signal \U409_TICK.TICK603_10\ : std_logic;
signal \U409_TICK.TICK603_9\ : std_logic;
signal \U409_TICK.TICK603_14\ : std_logic;
signal \TICK60_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \U409_TICK.TICK503_8\ : std_logic;
signal \U409_TICK.TICK503_11_cascade_\ : std_logic;
signal \U409_TICK.TICK503_14_cascade_\ : std_logic;
signal \TICK50_c\ : std_logic;
signal \U409_TICK.TICK503_9_cascade_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_0\ : std_logic;
signal \bfn_17_5_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_2\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_1\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_3\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_2\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_4\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_3\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_5\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_5\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_4\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_6\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_6\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_5\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_6\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_8\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_7\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_8\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_9\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_9\ : std_logic;
signal \bfn_17_6_0_\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_10\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_9\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_10\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_12\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_13\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_13\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_12\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_14\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_13\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_15\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_15\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_14\ : std_logic;
signal \U409_TICK.un2_COUNTER50_1_cry_15\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_16\ : std_logic;
signal \U409_TICK.TICK503_14\ : std_logic;
signal \U409_TICK.TICK503_9\ : std_logic;
signal \U409_TICK.TICK503_10\ : std_logic;
signal \U409_TICK.COUNTER50_RNO_0Z0Z_11\ : std_logic;
signal \U409_TICK.COUNTER50Z0Z_11\ : std_logic;
signal \CLK6_c_g\ : std_logic;
signal \PCS0_c\ : std_logic;
signal \SCS1_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z0\ : std_logic;
signal \PCS1_c\ : std_logic;
signal \U409_ADDRESS_DECODE.CSZ0Z1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \SCS0_c\ : std_logic;
signal \XCLK_ENn_c\ : std_logic;
signal \XCLK_c\ : std_logic;
signal \CLK28_IN_c_g\ : std_logic;
signal \AGNUS_CLK_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \CLK40_IN_wire\ : std_logic;
signal \CLK28_IN_wire\ : std_logic;
signal \CLK6_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(31 downto 1);
signal \TT_wire\ : std_logic_vector(1 downto 0);
signal \ROM_DELAY_wire\ : std_logic_vector(1 downto 0);
signal \CPUCONFn_wire\ : std_logic;
signal \RTC_ENn_wire\ : std_logic;
signal \SPIO_J_wire\ : std_logic;
signal \PPIO_wire\ : std_logic;
signal \TM_wire\ : std_logic_vector(2 downto 0);
signal \PPIO_J_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \ROMENn_wire\ : std_logic;
signal \TBIn_wire\ : std_logic;
signal \AUTOBOOT_wire\ : std_logic;
signal \F_READn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \PORTSIZE_wire\ : std_logic;
signal \F_ENn_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \SCS1_wire\ : std_logic;
signal \AGNUS_CLK_wire\ : std_logic;
signal \CIACS0n_wire\ : std_logic;
signal \TICK50_wire\ : std_logic;
signal \BREG_ENn_wire\ : std_logic;
signal \F_BANK_wire\ : std_logic_vector(1 downto 0);
signal \XCLK_ENn_wire\ : std_logic;
signal \TICK60_wire\ : std_logic;
signal \ATA_ENn_wire\ : std_logic;
signal \CIACS1n_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \PCS0_wire\ : std_logic;
signal \PCIAT_wire\ : std_logic_vector(1 downto 0);
signal \CLK_CIA_wire\ : std_logic;
signal \PCS1_wire\ : std_logic;
signal \BUFENn_wire\ : std_logic;
signal \F_WRITEn_wire\ : std_logic;
signal \SCS0_wire\ : std_logic;
signal \BPRO_ENn_wire\ : std_logic;
signal \XCLK_wire\ : std_logic;
signal \F_WPn_wire\ : std_logic;
signal \OVL_wire\ : std_logic;
signal \TCIn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \CONFIGENn_wire\ : std_logic;
signal \SPIO_wire\ : std_logic;
signal \F_RSTn_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    \CLK40_IN_wire\ <= CLK40_IN;
    \CLK28_IN_wire\ <= CLK28_IN;
    \CLK6_wire\ <= CLK6;
    \A_wire\ <= A;
    \TT_wire\ <= TT;
    \ROM_DELAY_wire\ <= ROM_DELAY;
    \CPUCONFn_wire\ <= CPUCONFn;
    RTC_ENn <= \RTC_ENn_wire\;
    \SPIO_J_wire\ <= SPIO_J;
    PPIO <= \PPIO_wire\;
    \TM_wire\ <= TM;
    \PPIO_J_wire\ <= PPIO_J;
    RAMSPACEn <= \RAMSPACEn_wire\;
    ROMENn <= \ROMENn_wire\;
    TBIn <= \TBIn_wire\;
    \AUTOBOOT_wire\ <= AUTOBOOT;
    F_READn <= \F_READn_wire\;
    \TSn_wire\ <= TSn;
    PORTSIZE <= \PORTSIZE_wire\;
    F_ENn <= \F_ENn_wire\;
    \RESETn_wire\ <= RESETn;
    SCS1 <= \SCS1_wire\;
    AGNUS_CLK <= \AGNUS_CLK_wire\;
    CIACS0n <= \CIACS0n_wire\;
    TICK50 <= \TICK50_wire\;
    BREG_ENn <= \BREG_ENn_wire\;
    F_BANK <= \F_BANK_wire\;
    \XCLK_ENn_wire\ <= XCLK_ENn;
    TICK60 <= \TICK60_wire\;
    ATA_ENn <= \ATA_ENn_wire\;
    CIACS1n <= \CIACS1n_wire\;
    REGSPACEn <= \REGSPACEn_wire\;
    PCS0 <= \PCS0_wire\;
    PCIAT <= \PCIAT_wire\;
    CLK_CIA <= \CLK_CIA_wire\;
    PCS1 <= \PCS1_wire\;
    BUFENn <= \BUFENn_wire\;
    F_WRITEn <= \F_WRITEn_wire\;
    SCS0 <= \SCS0_wire\;
    BPRO_ENn <= \BPRO_ENn_wire\;
    \XCLK_wire\ <= XCLK;
    F_WPn <= \F_WPn_wire\;
    \OVL_wire\ <= OVL;
    TCIn <= \TCIn_wire\;
    \RnW_wire\ <= RnW;
    CONFIGENn <= \CONFIGENn_wire\;
    SPIO <= \SPIO_wire\;
    F_RSTn <= \F_RSTn_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0001111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__8638\,
            RESETB => \N__11981\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => \CLK80_OUT\
        );

    \CLK40_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13651\,
            GLOBALBUFFEROUTPUT => \CLK40_IN_c_g\
        );

    \CLK40_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13653\,
            DIN => \N__13652\,
            DOUT => \N__13651\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13653\,
            PADOUT => \N__13652\,
            PADIN => \N__13651\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK28_IN_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13641\,
            GLOBALBUFFEROUTPUT => \CLK28_IN_c_g\
        );

    \CLK28_IN_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13643\,
            DIN => \N__13642\,
            DOUT => \N__13641\,
            PACKAGEPIN => \CLK28_IN_wire\
        );

    \CLK28_IN_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13643\,
            PADOUT => \N__13642\,
            PADIN => \N__13641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK6_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13631\,
            GLOBALBUFFEROUTPUT => \CLK6_c_g\
        );

    \CLK6_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13633\,
            DIN => \N__13632\,
            DOUT => \N__13631\,
            PACKAGEPIN => \CLK6_wire\
        );

    \CLK6_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13633\,
            PADOUT => \N__13632\,
            PADIN => \N__13631\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13622\,
            DIN => \N__13621\,
            DOUT => \N__13620\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13622\,
            PADOUT => \N__13621\,
            PADIN => \N__13620\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13613\,
            DIN => \N__13612\,
            DOUT => \N__13611\,
            PACKAGEPIN => \TT_wire\(0)
        );

    \TT_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13613\,
            PADOUT => \N__13612\,
            PADIN => \N__13611\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROM_DELAY_ibuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13604\,
            DIN => \N__13603\,
            DOUT => \N__13602\,
            PACKAGEPIN => \ROM_DELAY_wire\(1)
        );

    \ROM_DELAY_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13604\,
            PADOUT => \N__13603\,
            PADIN => \N__13602\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ROM_DELAY_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13595\,
            DIN => \N__13594\,
            DOUT => \N__13593\,
            PACKAGEPIN => D(7)
        );

    \D_iobuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13595\,
            PADOUT => \N__13594\,
            PADIN => \N__13593\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5236\,
            DIN0 => \D_in_7\,
            DOUT0 => \N__5836\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13586\,
            DIN => \N__13585\,
            DOUT => \N__13584\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13586\,
            PADOUT => \N__13585\,
            PADIN => \N__13584\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CPUCONFn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13577\,
            DIN => \N__13576\,
            DOUT => \N__13575\,
            PACKAGEPIN => \CPUCONFn_wire\
        );

    \CPUCONFn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13577\,
            PADOUT => \N__13576\,
            PADIN => \N__13575\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CPUCONFn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RTC_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13568\,
            DIN => \N__13567\,
            DOUT => \N__13566\,
            PACKAGEPIN => \RTC_ENn_wire\
        );

    \RTC_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13568\,
            PADOUT => \N__13567\,
            PADIN => \N__13566\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13559\,
            DIN => \N__13558\,
            DOUT => \N__13557\,
            PACKAGEPIN => \A_wire\(24)
        );

    \A_ibuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13559\,
            PADOUT => \N__13558\,
            PADIN => \N__13557\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_24\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13550\,
            DIN => \N__13549\,
            DOUT => \N__13548\,
            PACKAGEPIN => \SPIO_J_wire\
        );

    \SPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13550\,
            PADOUT => \N__13549\,
            PADIN => \N__13548\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13541\,
            DIN => \N__13540\,
            DOUT => \N__13539\,
            PACKAGEPIN => D(4)
        );

    \D_iobuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13541\,
            PADOUT => \N__13540\,
            PADIN => \N__13539\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5221\,
            DIN0 => \D_in_4\,
            DOUT0 => \N__6367\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13532\,
            DIN => \N__13531\,
            DOUT => \N__13530\,
            PACKAGEPIN => \PPIO_wire\
        );

    \PPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13532\,
            PADOUT => \N__13531\,
            PADIN => \N__13530\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4798\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13523\,
            DIN => \N__13522\,
            DOUT => \N__13521\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13523\,
            PADOUT => \N__13522\,
            PADIN => \N__13521\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13514\,
            DIN => \N__13513\,
            DOUT => \N__13512\,
            PACKAGEPIN => \TM_wire\(1)
        );

    \TM_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13514\,
            PADOUT => \N__13513\,
            PADIN => \N__13512\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13505\,
            DIN => \N__13504\,
            DOUT => \N__13503\,
            PACKAGEPIN => \A_wire\(21)
        );

    \A_ibuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13505\,
            PADOUT => \N__13504\,
            PADIN => \N__13503\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_21\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PPIO_J_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13496\,
            DIN => \N__13495\,
            DOUT => \N__13494\,
            PACKAGEPIN => \PPIO_J_wire\
        );

    \PPIO_J_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13496\,
            PADOUT => \N__13495\,
            PADIN => \N__13494\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \PPIO_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13487\,
            DIN => \N__13486\,
            DOUT => \N__13485\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13487\,
            PADOUT => \N__13486\,
            PADIN => \N__13485\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13478\,
            DIN => \N__13477\,
            DOUT => \N__13476\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13478\,
            PADOUT => \N__13477\,
            PADIN => \N__13476\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13469\,
            DIN => \N__13468\,
            DOUT => \N__13467\,
            PACKAGEPIN => \ROMENn_wire\
        );

    \ROMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13469\,
            PADOUT => \N__13468\,
            PADIN => \N__13467\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10291\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TBIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13460\,
            DIN => \N__13459\,
            DOUT => \N__13458\,
            PACKAGEPIN => \TBIn_wire\
        );

    \TBIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13460\,
            PADOUT => \N__13459\,
            PADIN => \N__13458\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9607\,
            DIN0 => OPEN,
            DOUT0 => \N__9498\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AUTOBOOT_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13451\,
            DIN => \N__13450\,
            DOUT => \N__13449\,
            PACKAGEPIN => \AUTOBOOT_wire\
        );

    \AUTOBOOT_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13451\,
            PADOUT => \N__13450\,
            PADIN => \N__13449\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AUTOBOOT_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_READn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13442\,
            DIN => \N__13441\,
            DOUT => \N__13440\,
            PACKAGEPIN => \F_READn_wire\
        );

    \F_READn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13442\,
            PADOUT => \N__13441\,
            PADIN => \N__13440\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12001\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13433\,
            DIN => \N__13432\,
            DOUT => \N__13431\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13433\,
            PADOUT => \N__13432\,
            PADIN => \N__13431\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PORTSIZE_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13424\,
            DIN => \N__13423\,
            DOUT => \N__13422\,
            PACKAGEPIN => \PORTSIZE_wire\
        );

    \PORTSIZE_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13424\,
            PADOUT => \N__13423\,
            PADIN => \N__13422\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5776\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13415\,
            DIN => \N__13414\,
            DOUT => \N__13413\,
            PACKAGEPIN => \F_ENn_wire\
        );

    \F_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13415\,
            PADOUT => \N__13414\,
            PADIN => \N__13413\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12000\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13406\,
            DIN => \N__13405\,
            DOUT => \N__13404\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13406\,
            PADOUT => \N__13405\,
            PADIN => \N__13404\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13397\,
            DIN => \N__13396\,
            DOUT => \N__13395\,
            PACKAGEPIN => \TM_wire\(2)
        );

    \TM_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13397\,
            PADOUT => \N__13396\,
            PADIN => \N__13395\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13388\,
            DIN => \N__13387\,
            DOUT => \N__13386\,
            PACKAGEPIN => \A_wire\(22)
        );

    \A_ibuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13388\,
            PADOUT => \N__13387\,
            PADIN => \N__13386\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_22\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13379\,
            DIN => \N__13378\,
            DOUT => \N__13377\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13379\,
            PADOUT => \N__13378\,
            PADIN => \N__13377\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13370\,
            DIN => \N__13369\,
            DOUT => \N__13368\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13370\,
            PADOUT => \N__13369\,
            PADIN => \N__13368\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13361\,
            DIN => \N__13360\,
            DOUT => \N__13359\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13361\,
            PADOUT => \N__13360\,
            PADIN => \N__13359\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ROM_DELAY_ibuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__13352\,
            DIN => \N__13351\,
            DOUT => \N__13350\,
            PACKAGEPIN => \ROM_DELAY_wire\(0)
        );

    \ROM_DELAY_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13352\,
            PADOUT => \N__13351\,
            PADIN => \N__13350\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \ROM_DELAY_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13343\,
            DIN => \N__13342\,
            DOUT => \N__13341\,
            PACKAGEPIN => \SCS1_wire\
        );

    \SCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13343\,
            PADOUT => \N__13342\,
            PADIN => \N__13341\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12553\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13334\,
            DIN => \N__13333\,
            DOUT => \N__13332\,
            PACKAGEPIN => \AGNUS_CLK_wire\
        );

    \AGNUS_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13334\,
            PADOUT => \N__13333\,
            PADIN => \N__13332\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12823\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13325\,
            DIN => \N__13324\,
            DOUT => \N__13323\,
            PACKAGEPIN => \A_wire\(25)
        );

    \A_ibuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13325\,
            PADOUT => \N__13324\,
            PADIN => \N__13323\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_25\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS0n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13316\,
            DIN => \N__13315\,
            DOUT => \N__13314\,
            PACKAGEPIN => \CIACS0n_wire\
        );

    \CIACS0n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13316\,
            PADOUT => \N__13315\,
            PADIN => \N__13314\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9124\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK50_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13307\,
            DIN => \N__13306\,
            DOUT => \N__13305\,
            PACKAGEPIN => \TICK50_wire\
        );

    \TICK50_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13307\,
            PADOUT => \N__13306\,
            PADIN => \N__13305\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12277\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13298\,
            DIN => \N__13297\,
            DOUT => \N__13296\,
            PACKAGEPIN => \A_wire\(28)
        );

    \A_ibuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13298\,
            PADOUT => \N__13297\,
            PADIN => \N__13296\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_28\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BREG_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13289\,
            DIN => \N__13288\,
            DOUT => \N__13287\,
            PACKAGEPIN => \BREG_ENn_wire\
        );

    \BREG_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13289\,
            PADOUT => \N__13288\,
            PADIN => \N__13287\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6565\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13280\,
            DIN => \N__13279\,
            DOUT => \N__13278\,
            PACKAGEPIN => D(5)
        );

    \D_iobuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13280\,
            PADOUT => \N__13279\,
            PADIN => \N__13278\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5231\,
            DIN0 => \D_in_5\,
            DOUT0 => \N__5404\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_BANK_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13271\,
            DIN => \N__13270\,
            DOUT => \N__13269\,
            PACKAGEPIN => \F_BANK_wire\(0)
        );

    \F_BANK_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13271\,
            PADOUT => \N__13270\,
            PADIN => \N__13269\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7144\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ENn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13262\,
            DIN => \N__13261\,
            DOUT => \N__13260\,
            PACKAGEPIN => \XCLK_ENn_wire\
        );

    \XCLK_ENn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13262\,
            PADOUT => \N__13261\,
            PADIN => \N__13260\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_ENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13253\,
            DIN => \N__13252\,
            DOUT => \N__13251\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13253\,
            PADOUT => \N__13252\,
            PADIN => \N__13251\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TICK60_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13244\,
            DIN => \N__13243\,
            DOUT => \N__13242\,
            PACKAGEPIN => \TICK60_wire\
        );

    \TICK60_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13244\,
            PADOUT => \N__13243\,
            PADIN => \N__13242\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12025\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13235\,
            DIN => \N__13234\,
            DOUT => \N__13233\,
            PACKAGEPIN => \A_wire\(26)
        );

    \A_ibuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13235\,
            PADOUT => \N__13234\,
            PADIN => \N__13233\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_26\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13226\,
            DIN => \N__13225\,
            DOUT => \N__13224\,
            PACKAGEPIN => \A_wire\(23)
        );

    \A_ibuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13226\,
            PADOUT => \N__13225\,
            PADIN => \N__13224\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_23\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13217\,
            DIN => \N__13216\,
            DOUT => \N__13215\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13217\,
            PADOUT => \N__13216\,
            PADIN => \N__13215\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ATA_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13208\,
            DIN => \N__13207\,
            DOUT => \N__13206\,
            PACKAGEPIN => \ATA_ENn_wire\
        );

    \ATA_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13208\,
            PADOUT => \N__13207\,
            PADIN => \N__13206\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8329\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13199\,
            DIN => \N__13198\,
            DOUT => \N__13197\,
            PACKAGEPIN => \A_wire\(31)
        );

    \A_ibuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13199\,
            PADOUT => \N__13198\,
            PADIN => \N__13197\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_31\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CIACS1n_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13190\,
            DIN => \N__13189\,
            DOUT => \N__13188\,
            PACKAGEPIN => \CIACS1n_wire\
        );

    \CIACS1n_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13190\,
            PADOUT => \N__13189\,
            PADIN => \N__13188\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13181\,
            DIN => \N__13180\,
            DOUT => \N__13179\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13181\,
            PADOUT => \N__13180\,
            PADIN => \N__13179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6652\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13172\,
            DIN => \N__13171\,
            DOUT => \N__13170\,
            PACKAGEPIN => \PCS0_wire\
        );

    \PCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13172\,
            PADOUT => \N__13171\,
            PADIN => \N__13170\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12571\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCIAT_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13163\,
            DIN => \N__13162\,
            DOUT => \N__13161\,
            PACKAGEPIN => \PCIAT_wire\(0)
        );

    \PCIAT_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13163\,
            PADOUT => \N__13162\,
            PADIN => \N__13161\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10465\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13154\,
            DIN => \N__13153\,
            DOUT => \N__13152\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13154\,
            PADOUT => \N__13153\,
            PADIN => \N__13152\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_CIA_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13145\,
            DIN => \N__13144\,
            DOUT => \N__13143\,
            PACKAGEPIN => \CLK_CIA_wire\
        );

    \CLK_CIA_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13145\,
            PADOUT => \N__13144\,
            PADIN => \N__13143\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13136\,
            DIN => \N__13135\,
            DOUT => \N__13134\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13136\,
            PADOUT => \N__13135\,
            PADIN => \N__13134\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCS1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13127\,
            DIN => \N__13126\,
            DOUT => \N__13125\,
            PACKAGEPIN => \PCS1_wire\
        );

    \PCS1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13127\,
            PADOUT => \N__13126\,
            PADIN => \N__13125\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12505\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_iobuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13118\,
            DIN => \N__13117\,
            DOUT => \N__13116\,
            PACKAGEPIN => TACKn
        );

    \TACKn_iobuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13118\,
            PADOUT => \N__13117\,
            PADIN => \N__13116\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9603\,
            DIN0 => \TACKn_in\,
            DOUT0 => \N__9491\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TT_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13109\,
            DIN => \N__13108\,
            DOUT => \N__13107\,
            PACKAGEPIN => \TT_wire\(1)
        );

    \TT_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13109\,
            PADOUT => \N__13108\,
            PADIN => \N__13107\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TT_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BUFENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13100\,
            DIN => \N__13099\,
            DOUT => \N__13098\,
            PACKAGEPIN => \BUFENn_wire\
        );

    \BUFENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13100\,
            PADOUT => \N__13099\,
            PADIN => \N__13098\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8377\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13091\,
            DIN => \N__13090\,
            DOUT => \N__13089\,
            PACKAGEPIN => \A_wire\(29)
        );

    \A_ibuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13091\,
            PADOUT => \N__13090\,
            PADIN => \N__13089\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_29\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \D_iobuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13082\,
            DIN => \N__13081\,
            DOUT => \N__13080\,
            PACKAGEPIN => D(6)
        );

    \D_iobuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__13082\,
            PADOUT => \N__13081\,
            PADIN => \N__13080\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__5232\,
            DIN0 => \D_in_6\,
            DOUT0 => \N__5422\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_BANK_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13073\,
            DIN => \N__13072\,
            DOUT => \N__13071\,
            PACKAGEPIN => \F_BANK_wire\(1)
        );

    \F_BANK_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13073\,
            PADOUT => \N__13072\,
            PADIN => \N__13071\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9049\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_WRITEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13064\,
            DIN => \N__13063\,
            DOUT => \N__13062\,
            PACKAGEPIN => \F_WRITEn_wire\
        );

    \F_WRITEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13064\,
            PADOUT => \N__13063\,
            PADIN => \N__13062\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11977\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13055\,
            DIN => \N__13054\,
            DOUT => \N__13053\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13055\,
            PADOUT => \N__13054\,
            PADIN => \N__13053\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13046\,
            DIN => \N__13045\,
            DOUT => \N__13044\,
            PACKAGEPIN => \A_wire\(27)
        );

    \A_ibuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13046\,
            PADOUT => \N__13045\,
            PADIN => \N__13044\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_27\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SCS0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13037\,
            DIN => \N__13036\,
            DOUT => \N__13035\,
            PACKAGEPIN => \SCS0_wire\
        );

    \SCS0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13037\,
            PADOUT => \N__13036\,
            PADIN => \N__13035\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12433\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BPRO_ENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13028\,
            DIN => \N__13027\,
            DOUT => \N__13026\,
            PACKAGEPIN => \BPRO_ENn_wire\
        );

    \BPRO_ENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13028\,
            PADOUT => \N__13027\,
            PADIN => \N__13026\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5143\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TM_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13019\,
            DIN => \N__13018\,
            DOUT => \N__13017\,
            PACKAGEPIN => \TM_wire\(0)
        );

    \TM_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13019\,
            PADOUT => \N__13018\,
            PADIN => \N__13017\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TM_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \XCLK_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13010\,
            DIN => \N__13009\,
            DOUT => \N__13008\,
            PACKAGEPIN => \XCLK_wire\
        );

    \XCLK_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13010\,
            PADOUT => \N__13009\,
            PADIN => \N__13008\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \XCLK_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13001\,
            DIN => \N__13000\,
            DOUT => \N__12999\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13001\,
            PADOUT => \N__13000\,
            PADIN => \N__12999\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_WPn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12992\,
            DIN => \N__12991\,
            DOUT => \N__12990\,
            PACKAGEPIN => \F_WPn_wire\
        );

    \F_WPn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12992\,
            PADOUT => \N__12991\,
            PADIN => \N__12990\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12983\,
            DIN => \N__12982\,
            DOUT => \N__12981\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12983\,
            PADOUT => \N__12982\,
            PADIN => \N__12981\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12974\,
            DIN => \N__12973\,
            DOUT => \N__12972\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12974\,
            PADOUT => \N__12973\,
            PADIN => \N__12972\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12965\,
            DIN => \N__12964\,
            DOUT => \N__12963\,
            PACKAGEPIN => \A_wire\(30)
        );

    \A_ibuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12965\,
            PADOUT => \N__12964\,
            PADIN => \N__12963\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_30\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \OVL_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12956\,
            DIN => \N__12955\,
            DOUT => \N__12954\,
            PACKAGEPIN => \OVL_wire\
        );

    \OVL_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12956\,
            PADOUT => \N__12955\,
            PADIN => \N__12954\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \OVL_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TCIn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12947\,
            DIN => \N__12946\,
            DOUT => \N__12945\,
            PACKAGEPIN => \TCIn_wire\
        );

    \TCIn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__12947\,
            PADOUT => \N__12946\,
            PADIN => \N__12945\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__9559\,
            DIN0 => OPEN,
            DOUT0 => \N__9499\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \PCIAT_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12938\,
            DIN => \N__12937\,
            DOUT => \N__12936\,
            PACKAGEPIN => \PCIAT_wire\(1)
        );

    \PCIAT_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12938\,
            PADOUT => \N__12937\,
            PADIN => \N__12936\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10555\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12929\,
            DIN => \N__12928\,
            DOUT => \N__12927\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12929\,
            PADOUT => \N__12928\,
            PADIN => \N__12927\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12920\,
            DIN => \N__12919\,
            DOUT => \N__12918\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12920\,
            PADOUT => \N__12919\,
            PADIN => \N__12918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CONFIGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12911\,
            DIN => \N__12910\,
            DOUT => \N__12909\,
            PACKAGEPIN => \CONFIGENn_wire\
        );

    \CONFIGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12911\,
            PADOUT => \N__12910\,
            PADIN => \N__12909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5194\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SPIO_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12902\,
            DIN => \N__12901\,
            DOUT => \N__12900\,
            PACKAGEPIN => \SPIO_wire\
        );

    \SPIO_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12902\,
            PADOUT => \N__12901\,
            PADIN => \N__12900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4777\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \F_RSTn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12893\,
            DIN => \N__12892\,
            DOUT => \N__12891\,
            PACKAGEPIN => \F_RSTn_wire\
        );

    \F_RSTn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12893\,
            PADOUT => \N__12892\,
            PADIN => \N__12891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11993\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3133\ : InMux
    port map (
            O => \N__12874\,
            I => \N__12871\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__12871\,
            I => \N__12868\
        );

    \I__3131\ : Span12Mux_v
    port map (
            O => \N__12868\,
            I => \N__12865\
        );

    \I__3130\ : Odrv12
    port map (
            O => \N__12865\,
            I => \XCLK_ENn_c\
        );

    \I__3129\ : InMux
    port map (
            O => \N__12862\,
            I => \N__12859\
        );

    \I__3128\ : LocalMux
    port map (
            O => \N__12859\,
            I => \N__12856\
        );

    \I__3127\ : Span4Mux_v
    port map (
            O => \N__12856\,
            I => \N__12853\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__12853\,
            I => \XCLK_c\
        );

    \I__3125\ : InMux
    port map (
            O => \N__12850\,
            I => \N__12847\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__12847\,
            I => \N__12840\
        );

    \I__3123\ : ClkMux
    port map (
            O => \N__12846\,
            I => \N__12829\
        );

    \I__3122\ : ClkMux
    port map (
            O => \N__12845\,
            I => \N__12829\
        );

    \I__3121\ : ClkMux
    port map (
            O => \N__12844\,
            I => \N__12829\
        );

    \I__3120\ : ClkMux
    port map (
            O => \N__12843\,
            I => \N__12829\
        );

    \I__3119\ : Glb2LocalMux
    port map (
            O => \N__12840\,
            I => \N__12829\
        );

    \I__3118\ : GlobalMux
    port map (
            O => \N__12829\,
            I => \N__12826\
        );

    \I__3117\ : gio2CtrlBuf
    port map (
            O => \N__12826\,
            I => \CLK28_IN_c_g\
        );

    \I__3116\ : IoInMux
    port map (
            O => \N__12823\,
            I => \N__12820\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__12820\,
            I => \N__12817\
        );

    \I__3114\ : Span4Mux_s3_h
    port map (
            O => \N__12817\,
            I => \N__12814\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__12814\,
            I => \AGNUS_CLK_c\
        );

    \I__3112\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12807\
        );

    \I__3111\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__12807\,
            I => \N__12801\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__12804\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__3108\ : Odrv4
    port map (
            O => \N__12801\,
            I => \U409_TICK.COUNTER50Z0Z_14\
        );

    \I__3107\ : InMux
    port map (
            O => \N__12796\,
            I => \N__12793\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__12793\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_14\
        );

    \I__3105\ : InMux
    port map (
            O => \N__12790\,
            I => \U409_TICK.un2_COUNTER50_1_cry_13\
        );

    \I__3104\ : InMux
    port map (
            O => \N__12787\,
            I => \N__12783\
        );

    \I__3103\ : InMux
    port map (
            O => \N__12786\,
            I => \N__12780\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__12783\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__12780\,
            I => \U409_TICK.COUNTER50Z0Z_15\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__12775\,
            I => \N__12772\
        );

    \I__3099\ : InMux
    port map (
            O => \N__12772\,
            I => \N__12769\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__12769\,
            I => \N__12766\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__12766\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_15\
        );

    \I__3096\ : InMux
    port map (
            O => \N__12763\,
            I => \U409_TICK.un2_COUNTER50_1_cry_14\
        );

    \I__3095\ : InMux
    port map (
            O => \N__12760\,
            I => \U409_TICK.un2_COUNTER50_1_cry_15\
        );

    \I__3094\ : InMux
    port map (
            O => \N__12757\,
            I => \N__12753\
        );

    \I__3093\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12750\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__12753\,
            I => \N__12747\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__12750\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__12747\,
            I => \U409_TICK.COUNTER50Z0Z_16\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__12742\,
            I => \N__12739\
        );

    \I__3088\ : InMux
    port map (
            O => \N__12739\,
            I => \N__12725\
        );

    \I__3087\ : InMux
    port map (
            O => \N__12738\,
            I => \N__12725\
        );

    \I__3086\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12725\
        );

    \I__3085\ : InMux
    port map (
            O => \N__12736\,
            I => \N__12716\
        );

    \I__3084\ : InMux
    port map (
            O => \N__12735\,
            I => \N__12716\
        );

    \I__3083\ : InMux
    port map (
            O => \N__12734\,
            I => \N__12716\
        );

    \I__3082\ : InMux
    port map (
            O => \N__12733\,
            I => \N__12716\
        );

    \I__3081\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12713\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__12725\,
            I => \U409_TICK.TICK503_14\
        );

    \I__3079\ : LocalMux
    port map (
            O => \N__12716\,
            I => \U409_TICK.TICK503_14\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__12713\,
            I => \U409_TICK.TICK503_14\
        );

    \I__3077\ : CascadeMux
    port map (
            O => \N__12706\,
            I => \N__12698\
        );

    \I__3076\ : InMux
    port map (
            O => \N__12705\,
            I => \N__12687\
        );

    \I__3075\ : InMux
    port map (
            O => \N__12704\,
            I => \N__12687\
        );

    \I__3074\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12687\
        );

    \I__3073\ : InMux
    port map (
            O => \N__12702\,
            I => \N__12687\
        );

    \I__3072\ : InMux
    port map (
            O => \N__12701\,
            I => \N__12684\
        );

    \I__3071\ : InMux
    port map (
            O => \N__12698\,
            I => \N__12677\
        );

    \I__3070\ : InMux
    port map (
            O => \N__12697\,
            I => \N__12677\
        );

    \I__3069\ : InMux
    port map (
            O => \N__12696\,
            I => \N__12677\
        );

    \I__3068\ : LocalMux
    port map (
            O => \N__12687\,
            I => \U409_TICK.TICK503_9\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__12684\,
            I => \U409_TICK.TICK503_9\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__12677\,
            I => \U409_TICK.TICK503_9\
        );

    \I__3065\ : CascadeMux
    port map (
            O => \N__12670\,
            I => \N__12665\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__12669\,
            I => \N__12657\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__12668\,
            I => \N__12654\
        );

    \I__3062\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12651\
        );

    \I__3061\ : InMux
    port map (
            O => \N__12664\,
            I => \N__12642\
        );

    \I__3060\ : InMux
    port map (
            O => \N__12663\,
            I => \N__12642\
        );

    \I__3059\ : InMux
    port map (
            O => \N__12662\,
            I => \N__12642\
        );

    \I__3058\ : InMux
    port map (
            O => \N__12661\,
            I => \N__12642\
        );

    \I__3057\ : InMux
    port map (
            O => \N__12660\,
            I => \N__12635\
        );

    \I__3056\ : InMux
    port map (
            O => \N__12657\,
            I => \N__12635\
        );

    \I__3055\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12635\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__12651\,
            I => \N__12632\
        );

    \I__3053\ : LocalMux
    port map (
            O => \N__12642\,
            I => \U409_TICK.TICK503_10\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__12635\,
            I => \U409_TICK.TICK503_10\
        );

    \I__3051\ : Odrv12
    port map (
            O => \N__12632\,
            I => \U409_TICK.TICK503_10\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12625\,
            I => \N__12622\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__12622\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_11\
        );

    \I__3048\ : InMux
    port map (
            O => \N__12619\,
            I => \N__12615\
        );

    \I__3047\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12612\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__12615\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__12612\,
            I => \U409_TICK.COUNTER50Z0Z_11\
        );

    \I__3044\ : ClkMux
    port map (
            O => \N__12607\,
            I => \N__12577\
        );

    \I__3043\ : ClkMux
    port map (
            O => \N__12606\,
            I => \N__12577\
        );

    \I__3042\ : ClkMux
    port map (
            O => \N__12605\,
            I => \N__12577\
        );

    \I__3041\ : ClkMux
    port map (
            O => \N__12604\,
            I => \N__12577\
        );

    \I__3040\ : ClkMux
    port map (
            O => \N__12603\,
            I => \N__12577\
        );

    \I__3039\ : ClkMux
    port map (
            O => \N__12602\,
            I => \N__12577\
        );

    \I__3038\ : ClkMux
    port map (
            O => \N__12601\,
            I => \N__12577\
        );

    \I__3037\ : ClkMux
    port map (
            O => \N__12600\,
            I => \N__12577\
        );

    \I__3036\ : ClkMux
    port map (
            O => \N__12599\,
            I => \N__12577\
        );

    \I__3035\ : ClkMux
    port map (
            O => \N__12598\,
            I => \N__12577\
        );

    \I__3034\ : GlobalMux
    port map (
            O => \N__12577\,
            I => \N__12574\
        );

    \I__3033\ : gio2CtrlBuf
    port map (
            O => \N__12574\,
            I => \CLK6_c_g\
        );

    \I__3032\ : IoInMux
    port map (
            O => \N__12571\,
            I => \N__12568\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__12568\,
            I => \N__12565\
        );

    \I__3030\ : IoSpan4Mux
    port map (
            O => \N__12565\,
            I => \N__12562\
        );

    \I__3029\ : Sp12to4
    port map (
            O => \N__12562\,
            I => \N__12559\
        );

    \I__3028\ : Span12Mux_s9_h
    port map (
            O => \N__12559\,
            I => \N__12556\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__12556\,
            I => \PCS0_c\
        );

    \I__3026\ : IoInMux
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__3024\ : IoSpan4Mux
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__3023\ : IoSpan4Mux
    port map (
            O => \N__12544\,
            I => \N__12541\
        );

    \I__3022\ : Span4Mux_s2_h
    port map (
            O => \N__12541\,
            I => \N__12538\
        );

    \I__3021\ : Span4Mux_h
    port map (
            O => \N__12538\,
            I => \N__12535\
        );

    \I__3020\ : Odrv4
    port map (
            O => \N__12535\,
            I => \SCS1_c\
        );

    \I__3019\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12529\
        );

    \I__3018\ : LocalMux
    port map (
            O => \N__12529\,
            I => \N__12525\
        );

    \I__3017\ : InMux
    port map (
            O => \N__12528\,
            I => \N__12522\
        );

    \I__3016\ : Span4Mux_v
    port map (
            O => \N__12525\,
            I => \N__12519\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__12522\,
            I => \N__12516\
        );

    \I__3014\ : Span4Mux_h
    port map (
            O => \N__12519\,
            I => \N__12513\
        );

    \I__3013\ : Span12Mux_s8_v
    port map (
            O => \N__12516\,
            I => \N__12510\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__12513\,
            I => \U409_ADDRESS_DECODE.CSZ0Z0\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__12510\,
            I => \U409_ADDRESS_DECODE.CSZ0Z0\
        );

    \I__3010\ : IoInMux
    port map (
            O => \N__12505\,
            I => \N__12502\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__12502\,
            I => \N__12499\
        );

    \I__3008\ : Span4Mux_s2_h
    port map (
            O => \N__12499\,
            I => \N__12496\
        );

    \I__3007\ : Sp12to4
    port map (
            O => \N__12496\,
            I => \N__12493\
        );

    \I__3006\ : Span12Mux_s7_v
    port map (
            O => \N__12493\,
            I => \N__12490\
        );

    \I__3005\ : Odrv12
    port map (
            O => \N__12490\,
            I => \PCS1_c\
        );

    \I__3004\ : InMux
    port map (
            O => \N__12487\,
            I => \N__12483\
        );

    \I__3003\ : InMux
    port map (
            O => \N__12486\,
            I => \N__12480\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__12483\,
            I => \N__12475\
        );

    \I__3001\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12475\
        );

    \I__3000\ : Odrv12
    port map (
            O => \N__12475\,
            I => \U409_ADDRESS_DECODE.CSZ0Z1\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12472\,
            I => \N__12466\
        );

    \I__2998\ : InMux
    port map (
            O => \N__12471\,
            I => \N__12463\
        );

    \I__2997\ : InMux
    port map (
            O => \N__12470\,
            I => \N__12460\
        );

    \I__2996\ : InMux
    port map (
            O => \N__12469\,
            I => \N__12457\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__12466\,
            I => \N__12452\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12463\,
            I => \N__12452\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__12460\,
            I => \N__12447\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__12457\,
            I => \N__12447\
        );

    \I__2991\ : Span4Mux_v
    port map (
            O => \N__12452\,
            I => \N__12444\
        );

    \I__2990\ : Span12Mux_v
    port map (
            O => \N__12447\,
            I => \N__12439\
        );

    \I__2989\ : Sp12to4
    port map (
            O => \N__12444\,
            I => \N__12439\
        );

    \I__2988\ : Span12Mux_h
    port map (
            O => \N__12439\,
            I => \N__12436\
        );

    \I__2987\ : Odrv12
    port map (
            O => \N__12436\,
            I => \A_c_14\
        );

    \I__2986\ : IoInMux
    port map (
            O => \N__12433\,
            I => \N__12430\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__12430\,
            I => \N__12427\
        );

    \I__2984\ : Span4Mux_s3_h
    port map (
            O => \N__12427\,
            I => \N__12424\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__12424\,
            I => \N__12421\
        );

    \I__2982\ : Span4Mux_h
    port map (
            O => \N__12421\,
            I => \N__12418\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__12418\,
            I => \SCS0_c\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__12415\,
            I => \N__12411\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__12414\,
            I => \N__12408\
        );

    \I__2978\ : InMux
    port map (
            O => \N__12411\,
            I => \N__12405\
        );

    \I__2977\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12402\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__12405\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__12402\,
            I => \U409_TICK.COUNTER50Z0Z_6\
        );

    \I__2974\ : InMux
    port map (
            O => \N__12397\,
            I => \N__12394\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__12394\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_6\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12391\,
            I => \U409_TICK.un2_COUNTER50_1_cry_5\
        );

    \I__2971\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12384\
        );

    \I__2970\ : InMux
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__2969\ : LocalMux
    port map (
            O => \N__12384\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__12381\,
            I => \U409_TICK.COUNTER50Z0Z_7\
        );

    \I__2967\ : InMux
    port map (
            O => \N__12376\,
            I => \U409_TICK.un2_COUNTER50_1_cry_6\
        );

    \I__2966\ : InMux
    port map (
            O => \N__12373\,
            I => \N__12369\
        );

    \I__2965\ : InMux
    port map (
            O => \N__12372\,
            I => \N__12366\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__12369\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2963\ : LocalMux
    port map (
            O => \N__12366\,
            I => \U409_TICK.COUNTER50Z0Z_8\
        );

    \I__2962\ : InMux
    port map (
            O => \N__12361\,
            I => \U409_TICK.un2_COUNTER50_1_cry_7\
        );

    \I__2961\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12354\
        );

    \I__2960\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__12354\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12351\,
            I => \U409_TICK.COUNTER50Z0Z_9\
        );

    \I__2957\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12343\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__12343\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_9\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12340\,
            I => \bfn_17_6_0_\
        );

    \I__2954\ : InMux
    port map (
            O => \N__12337\,
            I => \N__12334\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__12334\,
            I => \N__12330\
        );

    \I__2952\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12327\
        );

    \I__2951\ : Odrv4
    port map (
            O => \N__12330\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2950\ : LocalMux
    port map (
            O => \N__12327\,
            I => \U409_TICK.COUNTER50Z0Z_10\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12322\,
            I => \U409_TICK.un2_COUNTER50_1_cry_9\
        );

    \I__2948\ : InMux
    port map (
            O => \N__12319\,
            I => \U409_TICK.un2_COUNTER50_1_cry_10\
        );

    \I__2947\ : InMux
    port map (
            O => \N__12316\,
            I => \N__12313\
        );

    \I__2946\ : LocalMux
    port map (
            O => \N__12313\,
            I => \N__12309\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12312\,
            I => \N__12306\
        );

    \I__2944\ : Odrv4
    port map (
            O => \N__12309\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__12306\,
            I => \U409_TICK.COUNTER50Z0Z_12\
        );

    \I__2942\ : InMux
    port map (
            O => \N__12301\,
            I => \U409_TICK.un2_COUNTER50_1_cry_11\
        );

    \I__2941\ : InMux
    port map (
            O => \N__12298\,
            I => \N__12294\
        );

    \I__2940\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12291\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__12294\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__12291\,
            I => \U409_TICK.COUNTER50Z0Z_13\
        );

    \I__2937\ : InMux
    port map (
            O => \N__12286\,
            I => \N__12283\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__12283\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_13\
        );

    \I__2935\ : InMux
    port map (
            O => \N__12280\,
            I => \U409_TICK.un2_COUNTER50_1_cry_12\
        );

    \I__2934\ : IoInMux
    port map (
            O => \N__12277\,
            I => \N__12274\
        );

    \I__2933\ : LocalMux
    port map (
            O => \N__12274\,
            I => \N__12271\
        );

    \I__2932\ : Span4Mux_s1_v
    port map (
            O => \N__12271\,
            I => \N__12268\
        );

    \I__2931\ : Span4Mux_v
    port map (
            O => \N__12268\,
            I => \N__12265\
        );

    \I__2930\ : Span4Mux_v
    port map (
            O => \N__12265\,
            I => \N__12262\
        );

    \I__2929\ : Span4Mux_h
    port map (
            O => \N__12262\,
            I => \N__12258\
        );

    \I__2928\ : InMux
    port map (
            O => \N__12261\,
            I => \N__12255\
        );

    \I__2927\ : Odrv4
    port map (
            O => \N__12258\,
            I => \TICK50_c\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__12255\,
            I => \TICK50_c\
        );

    \I__2925\ : CascadeMux
    port map (
            O => \N__12250\,
            I => \U409_TICK.TICK503_9_cascade_\
        );

    \I__2924\ : InMux
    port map (
            O => \N__12247\,
            I => \N__12243\
        );

    \I__2923\ : InMux
    port map (
            O => \N__12246\,
            I => \N__12239\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__12243\,
            I => \N__12236\
        );

    \I__2921\ : InMux
    port map (
            O => \N__12242\,
            I => \N__12233\
        );

    \I__2920\ : LocalMux
    port map (
            O => \N__12239\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2919\ : Odrv4
    port map (
            O => \N__12236\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2918\ : LocalMux
    port map (
            O => \N__12233\,
            I => \U409_TICK.COUNTER50Z0Z_1\
        );

    \I__2917\ : InMux
    port map (
            O => \N__12226\,
            I => \N__12222\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__12225\,
            I => \N__12217\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__12222\,
            I => \N__12214\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12221\,
            I => \N__12209\
        );

    \I__2913\ : InMux
    port map (
            O => \N__12220\,
            I => \N__12209\
        );

    \I__2912\ : InMux
    port map (
            O => \N__12217\,
            I => \N__12206\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__12214\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__12209\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__12206\,
            I => \U409_TICK.COUNTER50Z0Z_0\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__12199\,
            I => \N__12196\
        );

    \I__2907\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12192\
        );

    \I__2906\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12189\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__12192\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__12189\,
            I => \U409_TICK.COUNTER50Z0Z_2\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12184\,
            I => \U409_TICK.un2_COUNTER50_1_cry_1\
        );

    \I__2902\ : InMux
    port map (
            O => \N__12181\,
            I => \N__12177\
        );

    \I__2901\ : InMux
    port map (
            O => \N__12180\,
            I => \N__12174\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__12177\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__12174\,
            I => \U409_TICK.COUNTER50Z0Z_3\
        );

    \I__2898\ : InMux
    port map (
            O => \N__12169\,
            I => \U409_TICK.un2_COUNTER50_1_cry_2\
        );

    \I__2897\ : CascadeMux
    port map (
            O => \N__12166\,
            I => \N__12163\
        );

    \I__2896\ : InMux
    port map (
            O => \N__12163\,
            I => \N__12159\
        );

    \I__2895\ : InMux
    port map (
            O => \N__12162\,
            I => \N__12156\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__12159\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__12156\,
            I => \U409_TICK.COUNTER50Z0Z_4\
        );

    \I__2892\ : InMux
    port map (
            O => \N__12151\,
            I => \U409_TICK.un2_COUNTER50_1_cry_3\
        );

    \I__2891\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12144\
        );

    \I__2890\ : InMux
    port map (
            O => \N__12147\,
            I => \N__12141\
        );

    \I__2889\ : LocalMux
    port map (
            O => \N__12144\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__12141\,
            I => \U409_TICK.COUNTER50Z0Z_5\
        );

    \I__2887\ : InMux
    port map (
            O => \N__12136\,
            I => \N__12133\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__12133\,
            I => \U409_TICK.COUNTER50_RNO_0Z0Z_5\
        );

    \I__2885\ : InMux
    port map (
            O => \N__12130\,
            I => \U409_TICK.un2_COUNTER50_1_cry_4\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__12127\,
            I => \U409_TICK.TICK503_10_cascade_\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__12124\,
            I => \N__12117\
        );

    \I__2882\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12112\
        );

    \I__2881\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12103\
        );

    \I__2880\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12103\
        );

    \I__2879\ : InMux
    port map (
            O => \N__12120\,
            I => \N__12103\
        );

    \I__2878\ : InMux
    port map (
            O => \N__12117\,
            I => \N__12103\
        );

    \I__2877\ : InMux
    port map (
            O => \N__12116\,
            I => \N__12098\
        );

    \I__2876\ : InMux
    port map (
            O => \N__12115\,
            I => \N__12098\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__12112\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__12103\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__12098\,
            I => \U409_TICK.TICK603_10\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12087\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__12090\,
            I => \N__12083\
        );

    \I__2870\ : InMux
    port map (
            O => \N__12087\,
            I => \N__12076\
        );

    \I__2869\ : InMux
    port map (
            O => \N__12086\,
            I => \N__12069\
        );

    \I__2868\ : InMux
    port map (
            O => \N__12083\,
            I => \N__12069\
        );

    \I__2867\ : InMux
    port map (
            O => \N__12082\,
            I => \N__12069\
        );

    \I__2866\ : InMux
    port map (
            O => \N__12081\,
            I => \N__12062\
        );

    \I__2865\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12062\
        );

    \I__2864\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12062\
        );

    \I__2863\ : LocalMux
    port map (
            O => \N__12076\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__12069\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__12062\,
            I => \U409_TICK.TICK603_9\
        );

    \I__2860\ : InMux
    port map (
            O => \N__12055\,
            I => \N__12046\
        );

    \I__2859\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12041\
        );

    \I__2858\ : InMux
    port map (
            O => \N__12053\,
            I => \N__12041\
        );

    \I__2857\ : InMux
    port map (
            O => \N__12052\,
            I => \N__12032\
        );

    \I__2856\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12032\
        );

    \I__2855\ : InMux
    port map (
            O => \N__12050\,
            I => \N__12032\
        );

    \I__2854\ : InMux
    port map (
            O => \N__12049\,
            I => \N__12032\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__12046\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__12041\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__12032\,
            I => \U409_TICK.TICK603_14\
        );

    \I__2850\ : IoInMux
    port map (
            O => \N__12025\,
            I => \N__12022\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__12022\,
            I => \N__12019\
        );

    \I__2848\ : Span4Mux_s3_v
    port map (
            O => \N__12019\,
            I => \N__12016\
        );

    \I__2847\ : Sp12to4
    port map (
            O => \N__12016\,
            I => \N__12013\
        );

    \I__2846\ : Span12Mux_h
    port map (
            O => \N__12013\,
            I => \N__12009\
        );

    \I__2845\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12006\
        );

    \I__2844\ : Odrv12
    port map (
            O => \N__12009\,
            I => \TICK60_c\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__12006\,
            I => \TICK60_c\
        );

    \I__2842\ : IoInMux
    port map (
            O => \N__12001\,
            I => \N__11997\
        );

    \I__2841\ : IoInMux
    port map (
            O => \N__12000\,
            I => \N__11994\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__11997\,
            I => \N__11988\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__2838\ : IoInMux
    port map (
            O => \N__11993\,
            I => \N__11985\
        );

    \I__2837\ : IoSpan4Mux
    port map (
            O => \N__11988\,
            I => \N__11982\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__11985\,
            I => \N__11978\
        );

    \I__2835\ : Span4Mux_s0_h
    port map (
            O => \N__11982\,
            I => \N__11974\
        );

    \I__2834\ : IoInMux
    port map (
            O => \N__11981\,
            I => \N__11971\
        );

    \I__2833\ : Span4Mux_s0_v
    port map (
            O => \N__11978\,
            I => \N__11968\
        );

    \I__2832\ : IoInMux
    port map (
            O => \N__11977\,
            I => \N__11965\
        );

    \I__2831\ : Sp12to4
    port map (
            O => \N__11974\,
            I => \N__11962\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__11971\,
            I => \N__11959\
        );

    \I__2829\ : Span4Mux_v
    port map (
            O => \N__11968\,
            I => \N__11956\
        );

    \I__2828\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11953\
        );

    \I__2827\ : Span12Mux_v
    port map (
            O => \N__11962\,
            I => \N__11948\
        );

    \I__2826\ : Span12Mux_s8_v
    port map (
            O => \N__11959\,
            I => \N__11948\
        );

    \I__2825\ : Span4Mux_v
    port map (
            O => \N__11956\,
            I => \N__11945\
        );

    \I__2824\ : Span12Mux_s8_v
    port map (
            O => \N__11953\,
            I => \N__11942\
        );

    \I__2823\ : Odrv12
    port map (
            O => \N__11948\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2822\ : Odrv4
    port map (
            O => \N__11945\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2821\ : Odrv12
    port map (
            O => \N__11942\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11935\,
            I => \N__11932\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__11932\,
            I => \U409_TICK.TICK503_8\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__11929\,
            I => \U409_TICK.TICK503_11_cascade_\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__11926\,
            I => \U409_TICK.TICK503_14_cascade_\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11923\,
            I => \N__11914\
        );

    \I__2815\ : InMux
    port map (
            O => \N__11922\,
            I => \N__11914\
        );

    \I__2814\ : InMux
    port map (
            O => \N__11921\,
            I => \N__11914\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__11914\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\
        );

    \I__2812\ : InMux
    port map (
            O => \N__11911\,
            I => \N__11905\
        );

    \I__2811\ : InMux
    port map (
            O => \N__11910\,
            I => \N__11898\
        );

    \I__2810\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11898\
        );

    \I__2809\ : InMux
    port map (
            O => \N__11908\,
            I => \N__11898\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11905\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__11898\,
            I => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\
        );

    \I__2806\ : InMux
    port map (
            O => \N__11893\,
            I => \N__11890\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__11890\,
            I => \U409_TRANSFER_ACK.N_3_0\
        );

    \I__2804\ : InMux
    port map (
            O => \N__11887\,
            I => \N__11884\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__11884\,
            I => \N__11880\
        );

    \I__2802\ : InMux
    port map (
            O => \N__11883\,
            I => \N__11877\
        );

    \I__2801\ : Span4Mux_v
    port map (
            O => \N__11880\,
            I => \N__11870\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__11877\,
            I => \N__11870\
        );

    \I__2799\ : InMux
    port map (
            O => \N__11876\,
            I => \N__11867\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11875\,
            I => \N__11864\
        );

    \I__2797\ : Span4Mux_v
    port map (
            O => \N__11870\,
            I => \N__11859\
        );

    \I__2796\ : LocalMux
    port map (
            O => \N__11867\,
            I => \N__11859\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__11864\,
            I => \N__11856\
        );

    \I__2794\ : Span4Mux_v
    port map (
            O => \N__11859\,
            I => \N__11843\
        );

    \I__2793\ : Span4Mux_v
    port map (
            O => \N__11856\,
            I => \N__11839\
        );

    \I__2792\ : InMux
    port map (
            O => \N__11855\,
            I => \N__11829\
        );

    \I__2791\ : InMux
    port map (
            O => \N__11854\,
            I => \N__11829\
        );

    \I__2790\ : InMux
    port map (
            O => \N__11853\,
            I => \N__11829\
        );

    \I__2789\ : InMux
    port map (
            O => \N__11852\,
            I => \N__11826\
        );

    \I__2788\ : InMux
    port map (
            O => \N__11851\,
            I => \N__11821\
        );

    \I__2787\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11821\
        );

    \I__2786\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11816\
        );

    \I__2785\ : InMux
    port map (
            O => \N__11848\,
            I => \N__11816\
        );

    \I__2784\ : InMux
    port map (
            O => \N__11847\,
            I => \N__11810\
        );

    \I__2783\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11810\
        );

    \I__2782\ : Span4Mux_h
    port map (
            O => \N__11843\,
            I => \N__11806\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11842\,
            I => \N__11803\
        );

    \I__2780\ : Span4Mux_h
    port map (
            O => \N__11839\,
            I => \N__11800\
        );

    \I__2779\ : InMux
    port map (
            O => \N__11838\,
            I => \N__11797\
        );

    \I__2778\ : InMux
    port map (
            O => \N__11837\,
            I => \N__11792\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__11836\,
            I => \N__11789\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__11829\,
            I => \N__11779\
        );

    \I__2775\ : LocalMux
    port map (
            O => \N__11826\,
            I => \N__11779\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11821\,
            I => \N__11779\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11779\
        );

    \I__2772\ : InMux
    port map (
            O => \N__11815\,
            I => \N__11776\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__11810\,
            I => \N__11772\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11809\,
            I => \N__11769\
        );

    \I__2769\ : Span4Mux_h
    port map (
            O => \N__11806\,
            I => \N__11764\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__11803\,
            I => \N__11764\
        );

    \I__2767\ : Span4Mux_h
    port map (
            O => \N__11800\,
            I => \N__11759\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__11797\,
            I => \N__11759\
        );

    \I__2765\ : InMux
    port map (
            O => \N__11796\,
            I => \N__11756\
        );

    \I__2764\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11753\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__11792\,
            I => \N__11750\
        );

    \I__2762\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11745\
        );

    \I__2761\ : InMux
    port map (
            O => \N__11788\,
            I => \N__11745\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__11779\,
            I => \N__11740\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__11776\,
            I => \N__11740\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__11775\,
            I => \N__11735\
        );

    \I__2757\ : Span4Mux_v
    port map (
            O => \N__11772\,
            I => \N__11732\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11728\
        );

    \I__2755\ : Span4Mux_v
    port map (
            O => \N__11764\,
            I => \N__11725\
        );

    \I__2754\ : Span4Mux_v
    port map (
            O => \N__11759\,
            I => \N__11722\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__11756\,
            I => \N__11719\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11716\
        );

    \I__2751\ : Span4Mux_h
    port map (
            O => \N__11750\,
            I => \N__11711\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__11745\,
            I => \N__11711\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__11740\,
            I => \N__11708\
        );

    \I__2748\ : InMux
    port map (
            O => \N__11739\,
            I => \N__11701\
        );

    \I__2747\ : InMux
    port map (
            O => \N__11738\,
            I => \N__11701\
        );

    \I__2746\ : InMux
    port map (
            O => \N__11735\,
            I => \N__11701\
        );

    \I__2745\ : Span4Mux_h
    port map (
            O => \N__11732\,
            I => \N__11698\
        );

    \I__2744\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11695\
        );

    \I__2743\ : Span12Mux_h
    port map (
            O => \N__11728\,
            I => \N__11692\
        );

    \I__2742\ : Sp12to4
    port map (
            O => \N__11725\,
            I => \N__11687\
        );

    \I__2741\ : Sp12to4
    port map (
            O => \N__11722\,
            I => \N__11687\
        );

    \I__2740\ : Span12Mux_v
    port map (
            O => \N__11719\,
            I => \N__11672\
        );

    \I__2739\ : Sp12to4
    port map (
            O => \N__11716\,
            I => \N__11672\
        );

    \I__2738\ : Sp12to4
    port map (
            O => \N__11711\,
            I => \N__11672\
        );

    \I__2737\ : Sp12to4
    port map (
            O => \N__11708\,
            I => \N__11672\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__11701\,
            I => \N__11672\
        );

    \I__2735\ : Sp12to4
    port map (
            O => \N__11698\,
            I => \N__11672\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__11695\,
            I => \N__11672\
        );

    \I__2733\ : Span12Mux_v
    port map (
            O => \N__11692\,
            I => \N__11669\
        );

    \I__2732\ : Span12Mux_h
    port map (
            O => \N__11687\,
            I => \N__11666\
        );

    \I__2731\ : Span12Mux_v
    port map (
            O => \N__11672\,
            I => \N__11663\
        );

    \I__2730\ : Span12Mux_h
    port map (
            O => \N__11669\,
            I => \N__11660\
        );

    \I__2729\ : Span12Mux_v
    port map (
            O => \N__11666\,
            I => \N__11655\
        );

    \I__2728\ : Span12Mux_h
    port map (
            O => \N__11663\,
            I => \N__11655\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11660\,
            I => \RESETn_c\
        );

    \I__2726\ : Odrv12
    port map (
            O => \N__11655\,
            I => \RESETn_c\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \N__11645\
        );

    \I__2724\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11640\
        );

    \I__2723\ : InMux
    port map (
            O => \N__11648\,
            I => \N__11640\
        );

    \I__2722\ : InMux
    port map (
            O => \N__11645\,
            I => \N__11637\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__11640\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__11637\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__11632\,
            I => \U409_TRANSFER_ACK.N_55_cascade_\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__11629\,
            I => \N__11622\
        );

    \I__2717\ : CascadeMux
    port map (
            O => \N__11628\,
            I => \N__11619\
        );

    \I__2716\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11616\
        );

    \I__2715\ : InMux
    port map (
            O => \N__11626\,
            I => \N__11607\
        );

    \I__2714\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11607\
        );

    \I__2713\ : InMux
    port map (
            O => \N__11622\,
            I => \N__11607\
        );

    \I__2712\ : InMux
    port map (
            O => \N__11619\,
            I => \N__11607\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__11616\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11607\,
            I => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\
        );

    \I__2709\ : InMux
    port map (
            O => \N__11602\,
            I => \N__11596\
        );

    \I__2708\ : InMux
    port map (
            O => \N__11601\,
            I => \N__11596\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__11596\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\
        );

    \I__2706\ : IoInMux
    port map (
            O => \N__11593\,
            I => \N__11590\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11587\
        );

    \I__2704\ : Span4Mux_s3_v
    port map (
            O => \N__11587\,
            I => \N__11583\
        );

    \I__2703\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__2702\ : Span4Mux_h
    port map (
            O => \N__11583\,
            I => \N__11577\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__11580\,
            I => \N__11574\
        );

    \I__2700\ : Span4Mux_h
    port map (
            O => \N__11577\,
            I => \N__11570\
        );

    \I__2699\ : Span4Mux_v
    port map (
            O => \N__11574\,
            I => \N__11567\
        );

    \I__2698\ : CascadeMux
    port map (
            O => \N__11573\,
            I => \N__11563\
        );

    \I__2697\ : Sp12to4
    port map (
            O => \N__11570\,
            I => \N__11560\
        );

    \I__2696\ : Span4Mux_h
    port map (
            O => \N__11567\,
            I => \N__11557\
        );

    \I__2695\ : InMux
    port map (
            O => \N__11566\,
            I => \N__11554\
        );

    \I__2694\ : InMux
    port map (
            O => \N__11563\,
            I => \N__11551\
        );

    \I__2693\ : Odrv12
    port map (
            O => \N__11560\,
            I => \CLK_CIA_c\
        );

    \I__2692\ : Odrv4
    port map (
            O => \N__11557\,
            I => \CLK_CIA_c\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__11554\,
            I => \CLK_CIA_c\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__11551\,
            I => \CLK_CIA_c\
        );

    \I__2689\ : InMux
    port map (
            O => \N__11542\,
            I => \N__11537\
        );

    \I__2688\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11532\
        );

    \I__2687\ : InMux
    port map (
            O => \N__11540\,
            I => \N__11532\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__11537\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2685\ : LocalMux
    port map (
            O => \N__11532\,
            I => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\
        );

    \I__2684\ : InMux
    port map (
            O => \N__11527\,
            I => \N__11524\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__11521\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11515\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11515\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__2678\ : InMux
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11506\,
            I => \N__11502\
        );

    \I__2676\ : InMux
    port map (
            O => \N__11505\,
            I => \N__11499\
        );

    \I__2675\ : Span4Mux_v
    port map (
            O => \N__11502\,
            I => \N__11494\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__11499\,
            I => \N__11491\
        );

    \I__2673\ : InMux
    port map (
            O => \N__11498\,
            I => \N__11488\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__11497\,
            I => \N__11485\
        );

    \I__2671\ : Span4Mux_h
    port map (
            O => \N__11494\,
            I => \N__11482\
        );

    \I__2670\ : Span4Mux_v
    port map (
            O => \N__11491\,
            I => \N__11479\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__11488\,
            I => \N__11476\
        );

    \I__2668\ : InMux
    port map (
            O => \N__11485\,
            I => \N__11473\
        );

    \I__2667\ : Odrv4
    port map (
            O => \N__11482\,
            I => \N_52_1\
        );

    \I__2666\ : Odrv4
    port map (
            O => \N__11479\,
            I => \N_52_1\
        );

    \I__2665\ : Odrv4
    port map (
            O => \N__11476\,
            I => \N_52_1\
        );

    \I__2664\ : LocalMux
    port map (
            O => \N__11473\,
            I => \N_52_1\
        );

    \I__2663\ : InMux
    port map (
            O => \N__11464\,
            I => \N__11460\
        );

    \I__2662\ : InMux
    port map (
            O => \N__11463\,
            I => \N__11455\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__11460\,
            I => \N__11452\
        );

    \I__2660\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11447\
        );

    \I__2659\ : InMux
    port map (
            O => \N__11458\,
            I => \N__11447\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__11455\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__2657\ : Odrv4
    port map (
            O => \N__11452\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11447\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\
        );

    \I__2655\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11437\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11431\
        );

    \I__2653\ : InMux
    port map (
            O => \N__11436\,
            I => \N__11426\
        );

    \I__2652\ : InMux
    port map (
            O => \N__11435\,
            I => \N__11421\
        );

    \I__2651\ : InMux
    port map (
            O => \N__11434\,
            I => \N__11421\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__11431\,
            I => \N__11417\
        );

    \I__2649\ : InMux
    port map (
            O => \N__11430\,
            I => \N__11412\
        );

    \I__2648\ : InMux
    port map (
            O => \N__11429\,
            I => \N__11412\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__11426\,
            I => \N__11407\
        );

    \I__2646\ : LocalMux
    port map (
            O => \N__11421\,
            I => \N__11407\
        );

    \I__2645\ : InMux
    port map (
            O => \N__11420\,
            I => \N__11404\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__11417\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11412\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__11407\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__11404\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\
        );

    \I__2640\ : SRMux
    port map (
            O => \N__11395\,
            I => \N__11353\
        );

    \I__2639\ : SRMux
    port map (
            O => \N__11394\,
            I => \N__11353\
        );

    \I__2638\ : SRMux
    port map (
            O => \N__11393\,
            I => \N__11353\
        );

    \I__2637\ : SRMux
    port map (
            O => \N__11392\,
            I => \N__11353\
        );

    \I__2636\ : SRMux
    port map (
            O => \N__11391\,
            I => \N__11353\
        );

    \I__2635\ : SRMux
    port map (
            O => \N__11390\,
            I => \N__11353\
        );

    \I__2634\ : SRMux
    port map (
            O => \N__11389\,
            I => \N__11353\
        );

    \I__2633\ : SRMux
    port map (
            O => \N__11388\,
            I => \N__11353\
        );

    \I__2632\ : SRMux
    port map (
            O => \N__11387\,
            I => \N__11353\
        );

    \I__2631\ : SRMux
    port map (
            O => \N__11386\,
            I => \N__11353\
        );

    \I__2630\ : SRMux
    port map (
            O => \N__11385\,
            I => \N__11353\
        );

    \I__2629\ : SRMux
    port map (
            O => \N__11384\,
            I => \N__11353\
        );

    \I__2628\ : SRMux
    port map (
            O => \N__11383\,
            I => \N__11353\
        );

    \I__2627\ : SRMux
    port map (
            O => \N__11382\,
            I => \N__11353\
        );

    \I__2626\ : GlobalMux
    port map (
            O => \N__11353\,
            I => \N__11350\
        );

    \I__2625\ : gio2CtrlBuf
    port map (
            O => \N__11350\,
            I => \RESETn_c_i_g\
        );

    \I__2624\ : InMux
    port map (
            O => \N__11347\,
            I => \N__11343\
        );

    \I__2623\ : InMux
    port map (
            O => \N__11346\,
            I => \N__11340\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__11343\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__11340\,
            I => \U409_TICK.COUNTER60Z0Z_12\
        );

    \I__2620\ : InMux
    port map (
            O => \N__11335\,
            I => \N__11331\
        );

    \I__2619\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11328\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__11331\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__11328\,
            I => \U409_TICK.COUNTER60Z0Z_2\
        );

    \I__2616\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11320\,
            I => \N__11316\
        );

    \I__2614\ : InMux
    port map (
            O => \N__11319\,
            I => \N__11312\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__11316\,
            I => \N__11309\
        );

    \I__2612\ : InMux
    port map (
            O => \N__11315\,
            I => \N__11306\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__11312\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2610\ : Odrv12
    port map (
            O => \N__11309\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__11306\,
            I => \U409_TICK.COUNTER60Z0Z_1\
        );

    \I__2608\ : InMux
    port map (
            O => \N__11299\,
            I => \N__11295\
        );

    \I__2607\ : InMux
    port map (
            O => \N__11298\,
            I => \N__11292\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__11295\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__11292\,
            I => \U409_TICK.COUNTER60Z0Z_16\
        );

    \I__2604\ : InMux
    port map (
            O => \N__11287\,
            I => \N__11284\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__11284\,
            I => \U409_TICK.TICK603_8\
        );

    \I__2602\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11277\
        );

    \I__2601\ : InMux
    port map (
            O => \N__11280\,
            I => \N__11274\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__11277\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__11274\,
            I => \U409_TICK.COUNTER60Z0Z_11\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__11269\,
            I => \U409_TICK.TICK603_11_cascade_\
        );

    \I__2597\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11262\
        );

    \I__2596\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11259\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__11262\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__11259\,
            I => \U409_TICK.COUNTER60Z0Z_3\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__11254\,
            I => \U409_TICK.TICK603_14_cascade_\
        );

    \I__2592\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11248\
        );

    \I__2591\ : LocalMux
    port map (
            O => \N__11248\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_14\
        );

    \I__2590\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11241\
        );

    \I__2589\ : InMux
    port map (
            O => \N__11244\,
            I => \N__11238\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__11241\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__11238\,
            I => \U409_TICK.COUNTER60Z0Z_14\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__11233\,
            I => \N__11230\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11230\,
            I => \N__11227\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__11227\,
            I => \N__11224\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__11224\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_15\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11221\,
            I => \N__11217\
        );

    \I__2581\ : InMux
    port map (
            O => \N__11220\,
            I => \N__11214\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__11217\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11214\,
            I => \U409_TICK.COUNTER60Z0Z_15\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__11209\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\
        );

    \I__2577\ : InMux
    port map (
            O => \N__11206\,
            I => \N__11199\
        );

    \I__2576\ : InMux
    port map (
            O => \N__11205\,
            I => \N__11196\
        );

    \I__2575\ : InMux
    port map (
            O => \N__11204\,
            I => \N__11191\
        );

    \I__2574\ : InMux
    port map (
            O => \N__11203\,
            I => \N__11191\
        );

    \I__2573\ : InMux
    port map (
            O => \N__11202\,
            I => \N__11188\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__11199\,
            I => \N__11184\
        );

    \I__2571\ : LocalMux
    port map (
            O => \N__11196\,
            I => \N__11176\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__11191\,
            I => \N__11166\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11188\,
            I => \N__11162\
        );

    \I__2568\ : ClkMux
    port map (
            O => \N__11187\,
            I => \N__11122\
        );

    \I__2567\ : Glb2LocalMux
    port map (
            O => \N__11184\,
            I => \N__11122\
        );

    \I__2566\ : ClkMux
    port map (
            O => \N__11183\,
            I => \N__11122\
        );

    \I__2565\ : ClkMux
    port map (
            O => \N__11182\,
            I => \N__11122\
        );

    \I__2564\ : ClkMux
    port map (
            O => \N__11181\,
            I => \N__11122\
        );

    \I__2563\ : ClkMux
    port map (
            O => \N__11180\,
            I => \N__11122\
        );

    \I__2562\ : ClkMux
    port map (
            O => \N__11179\,
            I => \N__11122\
        );

    \I__2561\ : Glb2LocalMux
    port map (
            O => \N__11176\,
            I => \N__11122\
        );

    \I__2560\ : ClkMux
    port map (
            O => \N__11175\,
            I => \N__11122\
        );

    \I__2559\ : ClkMux
    port map (
            O => \N__11174\,
            I => \N__11122\
        );

    \I__2558\ : ClkMux
    port map (
            O => \N__11173\,
            I => \N__11122\
        );

    \I__2557\ : ClkMux
    port map (
            O => \N__11172\,
            I => \N__11122\
        );

    \I__2556\ : ClkMux
    port map (
            O => \N__11171\,
            I => \N__11122\
        );

    \I__2555\ : ClkMux
    port map (
            O => \N__11170\,
            I => \N__11122\
        );

    \I__2554\ : ClkMux
    port map (
            O => \N__11169\,
            I => \N__11122\
        );

    \I__2553\ : Glb2LocalMux
    port map (
            O => \N__11166\,
            I => \N__11122\
        );

    \I__2552\ : ClkMux
    port map (
            O => \N__11165\,
            I => \N__11122\
        );

    \I__2551\ : Glb2LocalMux
    port map (
            O => \N__11162\,
            I => \N__11122\
        );

    \I__2550\ : ClkMux
    port map (
            O => \N__11161\,
            I => \N__11122\
        );

    \I__2549\ : GlobalMux
    port map (
            O => \N__11122\,
            I => \N__11119\
        );

    \I__2548\ : gio2CtrlBuf
    port map (
            O => \N__11119\,
            I => \CLK40_IN_c_g\
        );

    \I__2547\ : InMux
    port map (
            O => \N__11116\,
            I => \N__11112\
        );

    \I__2546\ : InMux
    port map (
            O => \N__11115\,
            I => \N__11109\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__11112\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__11109\,
            I => \U409_TRANSFER_ACK.N_17_mux\
        );

    \I__2543\ : CascadeMux
    port map (
            O => \N__11104\,
            I => \U409_TRANSFER_ACK.N_3_0_cascade_\
        );

    \I__2542\ : InMux
    port map (
            O => \N__11101\,
            I => \N__11098\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__11098\,
            I => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\
        );

    \I__2540\ : CascadeMux
    port map (
            O => \N__11095\,
            I => \N__11092\
        );

    \I__2539\ : InMux
    port map (
            O => \N__11092\,
            I => \N__11089\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__11089\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_8\
        );

    \I__2537\ : InMux
    port map (
            O => \N__11086\,
            I => \N__11082\
        );

    \I__2536\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11079\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__11082\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__11079\,
            I => \U409_TICK.COUNTER60Z0Z_5\
        );

    \I__2533\ : InMux
    port map (
            O => \N__11074\,
            I => \N__11071\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__11071\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_4\
        );

    \I__2531\ : InMux
    port map (
            O => \N__11068\,
            I => \N__11064\
        );

    \I__2530\ : InMux
    port map (
            O => \N__11067\,
            I => \N__11061\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__11064\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__11061\,
            I => \U409_TICK.COUNTER60Z0Z_4\
        );

    \I__2527\ : InMux
    port map (
            O => \N__11056\,
            I => \N__11052\
        );

    \I__2526\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11049\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__11052\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__11049\,
            I => \U409_TICK.COUNTER60Z0Z_9\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__11044\,
            I => \N__11040\
        );

    \I__2522\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11037\
        );

    \I__2521\ : InMux
    port map (
            O => \N__11040\,
            I => \N__11034\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__11037\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__11034\,
            I => \U409_TICK.COUNTER60Z0Z_8\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__11029\,
            I => \U409_TICK.TICK603_9_cascade_\
        );

    \I__2517\ : InMux
    port map (
            O => \N__11026\,
            I => \N__11023\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__11023\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_6\
        );

    \I__2515\ : CascadeMux
    port map (
            O => \N__11020\,
            I => \N__11017\
        );

    \I__2514\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11013\
        );

    \I__2513\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11010\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__11013\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__11010\,
            I => \U409_TICK.COUNTER60Z0Z_6\
        );

    \I__2510\ : InMux
    port map (
            O => \N__11005\,
            I => \N__11001\
        );

    \I__2509\ : InMux
    port map (
            O => \N__11004\,
            I => \N__10998\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__11001\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10998\,
            I => \U409_TICK.COUNTER60Z0Z_13\
        );

    \I__2506\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10989\
        );

    \I__2505\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10986\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__10989\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10986\,
            I => \U409_TICK.COUNTER60Z0Z_10\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__2501\ : InMux
    port map (
            O => \N__10978\,
            I => \N__10974\
        );

    \I__2500\ : InMux
    port map (
            O => \N__10977\,
            I => \N__10971\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__10974\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10971\,
            I => \U409_TICK.COUNTER60Z0Z_7\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__10966\,
            I => \U409_TICK.TICK603_10_cascade_\
        );

    \I__2496\ : CascadeMux
    port map (
            O => \N__10963\,
            I => \N__10957\
        );

    \I__2495\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10954\
        );

    \I__2494\ : InMux
    port map (
            O => \N__10961\,
            I => \N__10949\
        );

    \I__2493\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10949\
        );

    \I__2492\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10946\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10954\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2490\ : LocalMux
    port map (
            O => \N__10949\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__10946\,
            I => \U409_TICK.COUNTER60Z0Z_0\
        );

    \I__2488\ : InMux
    port map (
            O => \N__10939\,
            I => \N__10935\
        );

    \I__2487\ : InMux
    port map (
            O => \N__10938\,
            I => \N__10932\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10935\,
            I => \N__10929\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10932\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__10929\,
            I => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\
        );

    \I__2483\ : InMux
    port map (
            O => \N__10924\,
            I => \N__10920\
        );

    \I__2482\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10917\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__10920\,
            I => \N__10914\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__10917\,
            I => \N__10911\
        );

    \I__2479\ : Span4Mux_v
    port map (
            O => \N__10914\,
            I => \N__10908\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__10911\,
            I => \N__10905\
        );

    \I__2477\ : Span4Mux_v
    port map (
            O => \N__10908\,
            I => \N__10901\
        );

    \I__2476\ : Sp12to4
    port map (
            O => \N__10905\,
            I => \N__10898\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10904\,
            I => \N__10895\
        );

    \I__2474\ : Odrv4
    port map (
            O => \N__10901\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2473\ : Odrv12
    port map (
            O => \N__10898\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__10895\,
            I => \U409_CIA.VMAZ0\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10888\,
            I => \N__10884\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__10887\,
            I => \N__10881\
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__10884\,
            I => \N__10878\
        );

    \I__2468\ : InMux
    port map (
            O => \N__10881\,
            I => \N__10875\
        );

    \I__2467\ : Span4Mux_h
    port map (
            O => \N__10878\,
            I => \N__10870\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10875\,
            I => \N__10870\
        );

    \I__2465\ : Odrv4
    port map (
            O => \N__10870\,
            I => \U409_TRANSFER_ACK.N_33\
        );

    \I__2464\ : InMux
    port map (
            O => \N__10867\,
            I => \N__10864\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__10864\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0\
        );

    \I__2462\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10855\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__10860\,
            I => \N__10852\
        );

    \I__2460\ : InMux
    port map (
            O => \N__10859\,
            I => \N__10845\
        );

    \I__2459\ : InMux
    port map (
            O => \N__10858\,
            I => \N__10842\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10855\,
            I => \N__10839\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10852\,
            I => \N__10834\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10851\,
            I => \N__10834\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10850\,
            I => \N__10829\
        );

    \I__2454\ : InMux
    port map (
            O => \N__10849\,
            I => \N__10829\
        );

    \I__2453\ : InMux
    port map (
            O => \N__10848\,
            I => \N__10826\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__10845\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10842\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__10839\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__10834\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__10829\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10826\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\
        );

    \I__2446\ : InMux
    port map (
            O => \N__10813\,
            I => \N__10809\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10812\,
            I => \N__10802\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__10809\,
            I => \N__10799\
        );

    \I__2443\ : CascadeMux
    port map (
            O => \N__10808\,
            I => \N__10796\
        );

    \I__2442\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10792\
        );

    \I__2441\ : InMux
    port map (
            O => \N__10806\,
            I => \N__10789\
        );

    \I__2440\ : InMux
    port map (
            O => \N__10805\,
            I => \N__10786\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__10802\,
            I => \N__10783\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__10799\,
            I => \N__10780\
        );

    \I__2437\ : InMux
    port map (
            O => \N__10796\,
            I => \N__10777\
        );

    \I__2436\ : InMux
    port map (
            O => \N__10795\,
            I => \N__10774\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__10792\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10789\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2433\ : LocalMux
    port map (
            O => \N__10786\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2432\ : Odrv4
    port map (
            O => \N__10783\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2431\ : Odrv4
    port map (
            O => \N__10780\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10777\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__10774\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\
        );

    \I__2428\ : InMux
    port map (
            O => \N__10759\,
            I => \N__10751\
        );

    \I__2427\ : InMux
    port map (
            O => \N__10758\,
            I => \N__10748\
        );

    \I__2426\ : InMux
    port map (
            O => \N__10757\,
            I => \N__10745\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10756\,
            I => \N__10742\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10755\,
            I => \N__10737\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10754\,
            I => \N__10737\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__10751\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10748\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__10745\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10742\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2418\ : LocalMux
    port map (
            O => \N__10737\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__10726\,
            I => \N__10723\
        );

    \I__2416\ : InMux
    port map (
            O => \N__10723\,
            I => \N__10720\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10720\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__10717\,
            I => \N__10712\
        );

    \I__2413\ : CascadeMux
    port map (
            O => \N__10716\,
            I => \N__10709\
        );

    \I__2412\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10704\
        );

    \I__2411\ : InMux
    port map (
            O => \N__10712\,
            I => \N__10701\
        );

    \I__2410\ : InMux
    port map (
            O => \N__10709\,
            I => \N__10698\
        );

    \I__2409\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10695\
        );

    \I__2408\ : InMux
    port map (
            O => \N__10707\,
            I => \N__10692\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__10704\,
            I => \N__10687\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10687\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10698\,
            I => \N__10682\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__10695\,
            I => \N__10682\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__10692\,
            I => \N__10679\
        );

    \I__2402\ : Span4Mux_v
    port map (
            O => \N__10687\,
            I => \N__10676\
        );

    \I__2401\ : Span4Mux_v
    port map (
            O => \N__10682\,
            I => \N__10673\
        );

    \I__2400\ : Span12Mux_v
    port map (
            O => \N__10679\,
            I => \N__10668\
        );

    \I__2399\ : Sp12to4
    port map (
            O => \N__10676\,
            I => \N__10668\
        );

    \I__2398\ : Sp12to4
    port map (
            O => \N__10673\,
            I => \N__10665\
        );

    \I__2397\ : Span12Mux_h
    port map (
            O => \N__10668\,
            I => \N__10662\
        );

    \I__2396\ : Span12Mux_h
    port map (
            O => \N__10665\,
            I => \N__10659\
        );

    \I__2395\ : Span12Mux_v
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__2394\ : Span12Mux_v
    port map (
            O => \N__10659\,
            I => \N__10653\
        );

    \I__2393\ : Odrv12
    port map (
            O => \N__10656\,
            I => \ROM_DELAY_c_0\
        );

    \I__2392\ : Odrv12
    port map (
            O => \N__10653\,
            I => \ROM_DELAY_c_0\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10648\,
            I => \N__10641\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10641\
        );

    \I__2389\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10638\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10641\,
            I => \N__10632\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10638\,
            I => \N__10632\
        );

    \I__2386\ : InMux
    port map (
            O => \N__10637\,
            I => \N__10629\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__10632\,
            I => \N__10623\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10629\,
            I => \N__10623\
        );

    \I__2383\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10620\
        );

    \I__2382\ : Span4Mux_h
    port map (
            O => \N__10623\,
            I => \N__10615\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10620\,
            I => \N__10615\
        );

    \I__2380\ : Sp12to4
    port map (
            O => \N__10615\,
            I => \N__10612\
        );

    \I__2379\ : Span12Mux_v
    port map (
            O => \N__10612\,
            I => \N__10609\
        );

    \I__2378\ : Span12Mux_h
    port map (
            O => \N__10609\,
            I => \N__10606\
        );

    \I__2377\ : Odrv12
    port map (
            O => \N__10606\,
            I => \ROM_DELAY_c_1\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__10603\,
            I => \N__10599\
        );

    \I__2375\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10596\
        );

    \I__2374\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10593\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10596\,
            I => \U409_TRANSFER_ACK.N_31_i\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10593\,
            I => \U409_TRANSFER_ACK.N_31_i\
        );

    \I__2371\ : InMux
    port map (
            O => \N__10588\,
            I => \N__10585\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__10585\,
            I => \U409_TICK.COUNTER60_RNO_0Z0Z_9\
        );

    \I__2369\ : InMux
    port map (
            O => \N__10582\,
            I => \U409_TICK.un3_COUNTER60_1_cry_7\
        );

    \I__2368\ : InMux
    port map (
            O => \N__10579\,
            I => \bfn_14_7_0_\
        );

    \I__2367\ : InMux
    port map (
            O => \N__10576\,
            I => \U409_TICK.un3_COUNTER60_1_cry_9\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10573\,
            I => \U409_TICK.un3_COUNTER60_1_cry_10\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10570\,
            I => \U409_TICK.un3_COUNTER60_1_cry_11\
        );

    \I__2364\ : InMux
    port map (
            O => \N__10567\,
            I => \U409_TICK.un3_COUNTER60_1_cry_12\
        );

    \I__2363\ : InMux
    port map (
            O => \N__10564\,
            I => \U409_TICK.un3_COUNTER60_1_cry_13\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10561\,
            I => \U409_TICK.un3_COUNTER60_1_cry_14\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10558\,
            I => \U409_TICK.un3_COUNTER60_1_cry_15\
        );

    \I__2360\ : IoInMux
    port map (
            O => \N__10555\,
            I => \N__10552\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10552\,
            I => \N__10549\
        );

    \I__2358\ : IoSpan4Mux
    port map (
            O => \N__10549\,
            I => \N__10546\
        );

    \I__2357\ : Sp12to4
    port map (
            O => \N__10546\,
            I => \N__10543\
        );

    \I__2356\ : Span12Mux_s7_v
    port map (
            O => \N__10543\,
            I => \N__10540\
        );

    \I__2355\ : Span12Mux_v
    port map (
            O => \N__10540\,
            I => \N__10537\
        );

    \I__2354\ : Odrv12
    port map (
            O => \N__10537\,
            I => \PCIAT_c_1\
        );

    \I__2353\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10530\
        );

    \I__2352\ : InMux
    port map (
            O => \N__10533\,
            I => \N__10527\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__10530\,
            I => \N__10522\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__10527\,
            I => \N__10522\
        );

    \I__2349\ : Span4Mux_v
    port map (
            O => \N__10522\,
            I => \N__10519\
        );

    \I__2348\ : Sp12to4
    port map (
            O => \N__10519\,
            I => \N__10516\
        );

    \I__2347\ : Span12Mux_h
    port map (
            O => \N__10516\,
            I => \N__10513\
        );

    \I__2346\ : Odrv12
    port map (
            O => \N__10513\,
            I => \TM_c_0\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10506\
        );

    \I__2344\ : InMux
    port map (
            O => \N__10509\,
            I => \N__10503\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10506\,
            I => \N__10498\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10503\,
            I => \N__10498\
        );

    \I__2341\ : Span4Mux_v
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__2340\ : Sp12to4
    port map (
            O => \N__10495\,
            I => \N__10492\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__10492\,
            I => \U409_ADDRESS_DECODE.N_58_mux\
        );

    \I__2338\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10486\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10486\,
            I => \N__10483\
        );

    \I__2336\ : Span4Mux_v
    port map (
            O => \N__10483\,
            I => \N__10479\
        );

    \I__2335\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10476\
        );

    \I__2334\ : Sp12to4
    port map (
            O => \N__10479\,
            I => \N__10471\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10476\,
            I => \N__10471\
        );

    \I__2332\ : Span12Mux_h
    port map (
            O => \N__10471\,
            I => \N__10468\
        );

    \I__2331\ : Odrv12
    port map (
            O => \N__10468\,
            I => \TM_c_1\
        );

    \I__2330\ : IoInMux
    port map (
            O => \N__10465\,
            I => \N__10462\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__10462\,
            I => \N__10459\
        );

    \I__2328\ : Span4Mux_s3_h
    port map (
            O => \N__10459\,
            I => \N__10456\
        );

    \I__2327\ : Sp12to4
    port map (
            O => \N__10456\,
            I => \N__10453\
        );

    \I__2326\ : Span12Mux_s11_v
    port map (
            O => \N__10453\,
            I => \N__10450\
        );

    \I__2325\ : Span12Mux_h
    port map (
            O => \N__10450\,
            I => \N__10447\
        );

    \I__2324\ : Odrv12
    port map (
            O => \N__10447\,
            I => \PCIAT_c_0\
        );

    \I__2323\ : InMux
    port map (
            O => \N__10444\,
            I => \U409_TICK.un3_COUNTER60_1_cry_1\
        );

    \I__2322\ : InMux
    port map (
            O => \N__10441\,
            I => \U409_TICK.un3_COUNTER60_1_cry_2\
        );

    \I__2321\ : InMux
    port map (
            O => \N__10438\,
            I => \U409_TICK.un3_COUNTER60_1_cry_3\
        );

    \I__2320\ : InMux
    port map (
            O => \N__10435\,
            I => \U409_TICK.un3_COUNTER60_1_cry_4\
        );

    \I__2319\ : InMux
    port map (
            O => \N__10432\,
            I => \U409_TICK.un3_COUNTER60_1_cry_5\
        );

    \I__2318\ : InMux
    port map (
            O => \N__10429\,
            I => \U409_TICK.un3_COUNTER60_1_cry_6\
        );

    \I__2317\ : InMux
    port map (
            O => \N__10426\,
            I => \N__10420\
        );

    \I__2316\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10420\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__10420\,
            I => \N__10417\
        );

    \I__2314\ : Span4Mux_v
    port map (
            O => \N__10417\,
            I => \N__10414\
        );

    \I__2313\ : Span4Mux_h
    port map (
            O => \N__10414\,
            I => \N__10411\
        );

    \I__2312\ : Odrv4
    port map (
            O => \N__10411\,
            I => \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__10408\,
            I => \N__10404\
        );

    \I__2310\ : CascadeMux
    port map (
            O => \N__10407\,
            I => \N__10401\
        );

    \I__2309\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10396\
        );

    \I__2308\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10396\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__10396\,
            I => \N__10391\
        );

    \I__2306\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10388\
        );

    \I__2305\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10385\
        );

    \I__2304\ : Span4Mux_v
    port map (
            O => \N__10391\,
            I => \N__10382\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__10388\,
            I => \N__10379\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10376\
        );

    \I__2301\ : Span4Mux_v
    port map (
            O => \N__10382\,
            I => \N__10373\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__10379\,
            I => \N__10370\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__10376\,
            I => \N__10367\
        );

    \I__2298\ : Sp12to4
    port map (
            O => \N__10373\,
            I => \N__10362\
        );

    \I__2297\ : Sp12to4
    port map (
            O => \N__10370\,
            I => \N__10362\
        );

    \I__2296\ : Span4Mux_h
    port map (
            O => \N__10367\,
            I => \N__10359\
        );

    \I__2295\ : Span12Mux_h
    port map (
            O => \N__10362\,
            I => \N__10354\
        );

    \I__2294\ : Sp12to4
    port map (
            O => \N__10359\,
            I => \N__10354\
        );

    \I__2293\ : Span12Mux_v
    port map (
            O => \N__10354\,
            I => \N__10351\
        );

    \I__2292\ : Odrv12
    port map (
            O => \N__10351\,
            I => \TSn_c\
        );

    \I__2291\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10344\
        );

    \I__2290\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10341\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__10344\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__10341\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\
        );

    \I__2287\ : CascadeMux
    port map (
            O => \N__10336\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_\
        );

    \I__2286\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10329\
        );

    \I__2285\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10326\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__10329\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__10326\,
            I => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\
        );

    \I__2282\ : InMux
    port map (
            O => \N__10321\,
            I => \N__10318\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__10318\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0\
        );

    \I__2280\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10311\
        );

    \I__2279\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10308\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__10311\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__10308\,
            I => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\
        );

    \I__2276\ : CascadeMux
    port map (
            O => \N__10303\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_\
        );

    \I__2275\ : CascadeMux
    port map (
            O => \N__10300\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\
        );

    \I__2274\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__10294\,
            I => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0\
        );

    \I__2272\ : IoInMux
    port map (
            O => \N__10291\,
            I => \N__10288\
        );

    \I__2271\ : LocalMux
    port map (
            O => \N__10288\,
            I => \N__10285\
        );

    \I__2270\ : IoSpan4Mux
    port map (
            O => \N__10285\,
            I => \N__10282\
        );

    \I__2269\ : Span4Mux_s2_v
    port map (
            O => \N__10282\,
            I => \N__10279\
        );

    \I__2268\ : Span4Mux_v
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__2267\ : Sp12to4
    port map (
            O => \N__10276\,
            I => \N__10272\
        );

    \I__2266\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10269\
        );

    \I__2265\ : Odrv12
    port map (
            O => \N__10272\,
            I => \ROMENn_c\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__10269\,
            I => \ROMENn_c\
        );

    \I__2263\ : InMux
    port map (
            O => \N__10264\,
            I => \N__10261\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__10261\,
            I => \U409_TRANSFER_ACK.N_42_i\
        );

    \I__2261\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10255\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10255\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\
        );

    \I__2259\ : InMux
    port map (
            O => \N__10252\,
            I => \N__10249\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__10249\,
            I => \N__10246\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__10246\,
            I => \N__10242\
        );

    \I__2256\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10239\
        );

    \I__2255\ : Odrv4
    port map (
            O => \N__10242\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_2\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__10239\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_2\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__10234\,
            I => \N__10231\
        );

    \I__2252\ : InMux
    port map (
            O => \N__10231\,
            I => \N__10228\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__10228\,
            I => \N__10225\
        );

    \I__2250\ : Odrv4
    port map (
            O => \N__10225\,
            I => \U409_ADDRESS_DECODE.N_61\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__10222\,
            I => \U409_TRANSFER_ACK.N_42_i_cascade_\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__10219\,
            I => \N__10215\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__10218\,
            I => \N__10210\
        );

    \I__2246\ : InMux
    port map (
            O => \N__10215\,
            I => \N__10206\
        );

    \I__2245\ : InMux
    port map (
            O => \N__10214\,
            I => \N__10203\
        );

    \I__2244\ : InMux
    port map (
            O => \N__10213\,
            I => \N__10198\
        );

    \I__2243\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10198\
        );

    \I__2242\ : InMux
    port map (
            O => \N__10209\,
            I => \N__10195\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10206\,
            I => \N__10191\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__10203\,
            I => \N__10187\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__10198\,
            I => \N__10184\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__10195\,
            I => \N__10181\
        );

    \I__2237\ : InMux
    port map (
            O => \N__10194\,
            I => \N__10178\
        );

    \I__2236\ : Span4Mux_v
    port map (
            O => \N__10191\,
            I => \N__10175\
        );

    \I__2235\ : InMux
    port map (
            O => \N__10190\,
            I => \N__10171\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__10187\,
            I => \N__10168\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__10184\,
            I => \N__10163\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__10181\,
            I => \N__10163\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__10178\,
            I => \N__10160\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__10175\,
            I => \N__10157\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10174\,
            I => \N__10154\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__10151\
        );

    \I__2227\ : Span4Mux_v
    port map (
            O => \N__10168\,
            I => \N__10148\
        );

    \I__2226\ : Span4Mux_h
    port map (
            O => \N__10163\,
            I => \N__10143\
        );

    \I__2225\ : Span4Mux_v
    port map (
            O => \N__10160\,
            I => \N__10143\
        );

    \I__2224\ : Span4Mux_h
    port map (
            O => \N__10157\,
            I => \N__10138\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__10154\,
            I => \N__10138\
        );

    \I__2222\ : Span12Mux_v
    port map (
            O => \N__10151\,
            I => \N__10135\
        );

    \I__2221\ : Sp12to4
    port map (
            O => \N__10148\,
            I => \N__10132\
        );

    \I__2220\ : Span4Mux_v
    port map (
            O => \N__10143\,
            I => \N__10129\
        );

    \I__2219\ : Sp12to4
    port map (
            O => \N__10138\,
            I => \N__10126\
        );

    \I__2218\ : Span12Mux_h
    port map (
            O => \N__10135\,
            I => \N__10123\
        );

    \I__2217\ : Span12Mux_h
    port map (
            O => \N__10132\,
            I => \N__10116\
        );

    \I__2216\ : Sp12to4
    port map (
            O => \N__10129\,
            I => \N__10116\
        );

    \I__2215\ : Span12Mux_v
    port map (
            O => \N__10126\,
            I => \N__10116\
        );

    \I__2214\ : Odrv12
    port map (
            O => \N__10123\,
            I => \A_c_23\
        );

    \I__2213\ : Odrv12
    port map (
            O => \N__10116\,
            I => \A_c_23\
        );

    \I__2212\ : InMux
    port map (
            O => \N__10111\,
            I => \N__10104\
        );

    \I__2211\ : InMux
    port map (
            O => \N__10110\,
            I => \N__10101\
        );

    \I__2210\ : InMux
    port map (
            O => \N__10109\,
            I => \N__10097\
        );

    \I__2209\ : InMux
    port map (
            O => \N__10108\,
            I => \N__10094\
        );

    \I__2208\ : InMux
    port map (
            O => \N__10107\,
            I => \N__10091\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10085\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__10101\,
            I => \N__10085\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10082\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__10097\,
            I => \N__10079\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__10094\,
            I => \N__10074\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10074\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10090\,
            I => \N__10071\
        );

    \I__2200\ : Span4Mux_v
    port map (
            O => \N__10085\,
            I => \N__10068\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__10082\,
            I => \N__10065\
        );

    \I__2198\ : Span4Mux_v
    port map (
            O => \N__10079\,
            I => \N__10062\
        );

    \I__2197\ : Span4Mux_v
    port map (
            O => \N__10074\,
            I => \N__10057\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__10071\,
            I => \N__10057\
        );

    \I__2195\ : Span4Mux_v
    port map (
            O => \N__10068\,
            I => \N__10054\
        );

    \I__2194\ : Span4Mux_v
    port map (
            O => \N__10065\,
            I => \N__10051\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__10062\,
            I => \N__10046\
        );

    \I__2192\ : Span4Mux_v
    port map (
            O => \N__10057\,
            I => \N__10046\
        );

    \I__2191\ : Span4Mux_h
    port map (
            O => \N__10054\,
            I => \N__10042\
        );

    \I__2190\ : Span4Mux_v
    port map (
            O => \N__10051\,
            I => \N__10037\
        );

    \I__2189\ : Span4Mux_h
    port map (
            O => \N__10046\,
            I => \N__10037\
        );

    \I__2188\ : InMux
    port map (
            O => \N__10045\,
            I => \N__10034\
        );

    \I__2187\ : Sp12to4
    port map (
            O => \N__10042\,
            I => \N__10027\
        );

    \I__2186\ : Sp12to4
    port map (
            O => \N__10037\,
            I => \N__10027\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__10034\,
            I => \N__10027\
        );

    \I__2184\ : Odrv12
    port map (
            O => \N__10027\,
            I => \A_c_20\
        );

    \I__2183\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10021\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__10021\,
            I => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__10018\,
            I => \N__10013\
        );

    \I__2180\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10006\
        );

    \I__2179\ : InMux
    port map (
            O => \N__10016\,
            I => \N__10002\
        );

    \I__2178\ : InMux
    port map (
            O => \N__10013\,
            I => \N__9999\
        );

    \I__2177\ : InMux
    port map (
            O => \N__10012\,
            I => \N__9996\
        );

    \I__2176\ : InMux
    port map (
            O => \N__10011\,
            I => \N__9993\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__10010\,
            I => \N__9990\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__10009\,
            I => \N__9987\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__10006\,
            I => \N__9984\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__10005\,
            I => \N__9981\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__10002\,
            I => \N__9978\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__9999\,
            I => \N__9975\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__9996\,
            I => \N__9969\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__9993\,
            I => \N__9969\
        );

    \I__2167\ : InMux
    port map (
            O => \N__9990\,
            I => \N__9966\
        );

    \I__2166\ : InMux
    port map (
            O => \N__9987\,
            I => \N__9963\
        );

    \I__2165\ : Span4Mux_v
    port map (
            O => \N__9984\,
            I => \N__9960\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9981\,
            I => \N__9957\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9978\,
            I => \N__9954\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9975\,
            I => \N__9951\
        );

    \I__2161\ : InMux
    port map (
            O => \N__9974\,
            I => \N__9948\
        );

    \I__2160\ : Span12Mux_v
    port map (
            O => \N__9969\,
            I => \N__9943\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__9966\,
            I => \N__9943\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9963\,
            I => \N__9930\
        );

    \I__2157\ : Sp12to4
    port map (
            O => \N__9960\,
            I => \N__9930\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9930\
        );

    \I__2155\ : Sp12to4
    port map (
            O => \N__9954\,
            I => \N__9930\
        );

    \I__2154\ : Sp12to4
    port map (
            O => \N__9951\,
            I => \N__9930\
        );

    \I__2153\ : LocalMux
    port map (
            O => \N__9948\,
            I => \N__9930\
        );

    \I__2152\ : Span12Mux_v
    port map (
            O => \N__9943\,
            I => \N__9927\
        );

    \I__2151\ : Span12Mux_h
    port map (
            O => \N__9930\,
            I => \N__9924\
        );

    \I__2150\ : Span12Mux_h
    port map (
            O => \N__9927\,
            I => \N__9919\
        );

    \I__2149\ : Span12Mux_v
    port map (
            O => \N__9924\,
            I => \N__9919\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__9919\,
            I => \A_c_19\
        );

    \I__2147\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9909\
        );

    \I__2146\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9906\
        );

    \I__2145\ : InMux
    port map (
            O => \N__9914\,
            I => \N__9903\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9900\
        );

    \I__2143\ : InMux
    port map (
            O => \N__9912\,
            I => \N__9896\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__9909\,
            I => \N__9892\
        );

    \I__2141\ : LocalMux
    port map (
            O => \N__9906\,
            I => \N__9889\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9903\,
            I => \N__9886\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__9900\,
            I => \N__9883\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9899\,
            I => \N__9880\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__9896\,
            I => \N__9877\
        );

    \I__2136\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9874\
        );

    \I__2135\ : Span4Mux_v
    port map (
            O => \N__9892\,
            I => \N__9871\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9889\,
            I => \N__9868\
        );

    \I__2133\ : Span4Mux_v
    port map (
            O => \N__9886\,
            I => \N__9864\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__9883\,
            I => \N__9861\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__9880\,
            I => \N__9854\
        );

    \I__2130\ : Span4Mux_h
    port map (
            O => \N__9877\,
            I => \N__9854\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9874\,
            I => \N__9854\
        );

    \I__2128\ : Span4Mux_v
    port map (
            O => \N__9871\,
            I => \N__9851\
        );

    \I__2127\ : Span4Mux_v
    port map (
            O => \N__9868\,
            I => \N__9848\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9845\
        );

    \I__2125\ : Sp12to4
    port map (
            O => \N__9864\,
            I => \N__9840\
        );

    \I__2124\ : Sp12to4
    port map (
            O => \N__9861\,
            I => \N__9840\
        );

    \I__2123\ : Sp12to4
    port map (
            O => \N__9854\,
            I => \N__9837\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__9851\,
            I => \N__9834\
        );

    \I__2121\ : Span4Mux_v
    port map (
            O => \N__9848\,
            I => \N__9831\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9845\,
            I => \N__9828\
        );

    \I__2119\ : Span12Mux_h
    port map (
            O => \N__9840\,
            I => \N__9825\
        );

    \I__2118\ : Span12Mux_v
    port map (
            O => \N__9837\,
            I => \N__9822\
        );

    \I__2117\ : Sp12to4
    port map (
            O => \N__9834\,
            I => \N__9819\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__9831\,
            I => \N__9816\
        );

    \I__2115\ : Sp12to4
    port map (
            O => \N__9828\,
            I => \N__9813\
        );

    \I__2114\ : Span12Mux_v
    port map (
            O => \N__9825\,
            I => \N__9808\
        );

    \I__2113\ : Span12Mux_h
    port map (
            O => \N__9822\,
            I => \N__9808\
        );

    \I__2112\ : Span12Mux_h
    port map (
            O => \N__9819\,
            I => \N__9801\
        );

    \I__2111\ : Sp12to4
    port map (
            O => \N__9816\,
            I => \N__9801\
        );

    \I__2110\ : Span12Mux_v
    port map (
            O => \N__9813\,
            I => \N__9801\
        );

    \I__2109\ : Odrv12
    port map (
            O => \N__9808\,
            I => \A_c_22\
        );

    \I__2108\ : Odrv12
    port map (
            O => \N__9801\,
            I => \A_c_22\
        );

    \I__2107\ : InMux
    port map (
            O => \N__9796\,
            I => \N__9792\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__9795\,
            I => \N__9789\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9786\
        );

    \I__2104\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9782\
        );

    \I__2103\ : Span4Mux_v
    port map (
            O => \N__9786\,
            I => \N__9779\
        );

    \I__2102\ : InMux
    port map (
            O => \N__9785\,
            I => \N__9776\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__9782\,
            I => \N__9769\
        );

    \I__2100\ : Sp12to4
    port map (
            O => \N__9779\,
            I => \N__9769\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9776\,
            I => \N__9769\
        );

    \I__2098\ : Span12Mux_v
    port map (
            O => \N__9769\,
            I => \N__9766\
        );

    \I__2097\ : Span12Mux_h
    port map (
            O => \N__9766\,
            I => \N__9763\
        );

    \I__2096\ : Odrv12
    port map (
            O => \N__9763\,
            I => \OVL_c\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__9760\,
            I => \N__9755\
        );

    \I__2094\ : InMux
    port map (
            O => \N__9759\,
            I => \N__9751\
        );

    \I__2093\ : InMux
    port map (
            O => \N__9758\,
            I => \N__9748\
        );

    \I__2092\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9745\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__9754\,
            I => \N__9741\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__9751\,
            I => \N__9733\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__9748\,
            I => \N__9733\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9745\,
            I => \N__9733\
        );

    \I__2087\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9730\
        );

    \I__2086\ : InMux
    port map (
            O => \N__9741\,
            I => \N__9725\
        );

    \I__2085\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9720\
        );

    \I__2084\ : Span4Mux_h
    port map (
            O => \N__9733\,
            I => \N__9715\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__9730\,
            I => \N__9715\
        );

    \I__2082\ : InMux
    port map (
            O => \N__9729\,
            I => \N__9712\
        );

    \I__2081\ : InMux
    port map (
            O => \N__9728\,
            I => \N__9709\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__9725\,
            I => \N__9705\
        );

    \I__2079\ : InMux
    port map (
            O => \N__9724\,
            I => \N__9702\
        );

    \I__2078\ : InMux
    port map (
            O => \N__9723\,
            I => \N__9699\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__9720\,
            I => \N__9695\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__9715\,
            I => \N__9690\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__9712\,
            I => \N__9690\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__9709\,
            I => \N__9687\
        );

    \I__2073\ : InMux
    port map (
            O => \N__9708\,
            I => \N__9684\
        );

    \I__2072\ : Span4Mux_v
    port map (
            O => \N__9705\,
            I => \N__9676\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__9702\,
            I => \N__9676\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__9699\,
            I => \N__9676\
        );

    \I__2069\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9673\
        );

    \I__2068\ : Span4Mux_h
    port map (
            O => \N__9695\,
            I => \N__9668\
        );

    \I__2067\ : Span4Mux_v
    port map (
            O => \N__9690\,
            I => \N__9668\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__9687\,
            I => \N__9665\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__9684\,
            I => \N__9662\
        );

    \I__2064\ : InMux
    port map (
            O => \N__9683\,
            I => \N__9659\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__9676\,
            I => \N__9656\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9673\,
            I => \N__9653\
        );

    \I__2061\ : Span4Mux_v
    port map (
            O => \N__9668\,
            I => \N__9646\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__9665\,
            I => \N__9646\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__9662\,
            I => \N__9646\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9659\,
            I => \N__9643\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__9656\,
            I => \N__9640\
        );

    \I__2056\ : Sp12to4
    port map (
            O => \N__9653\,
            I => \N__9637\
        );

    \I__2055\ : Span4Mux_h
    port map (
            O => \N__9646\,
            I => \N__9632\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__9643\,
            I => \N__9632\
        );

    \I__2053\ : Sp12to4
    port map (
            O => \N__9640\,
            I => \N__9625\
        );

    \I__2052\ : Span12Mux_v
    port map (
            O => \N__9637\,
            I => \N__9625\
        );

    \I__2051\ : Sp12to4
    port map (
            O => \N__9632\,
            I => \N__9625\
        );

    \I__2050\ : Odrv12
    port map (
            O => \N__9625\,
            I => \A_c_21\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9619\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9619\,
            I => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9616\,
            I => \N__9613\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__9613\,
            I => \N__9610\
        );

    \I__2045\ : Odrv12
    port map (
            O => \N__9610\,
            I => \ROMEN\
        );

    \I__2044\ : IoInMux
    port map (
            O => \N__9607\,
            I => \N__9604\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__9604\,
            I => \N__9600\
        );

    \I__2042\ : IoInMux
    port map (
            O => \N__9603\,
            I => \N__9597\
        );

    \I__2041\ : Span12Mux_s5_v
    port map (
            O => \N__9600\,
            I => \N__9594\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__9597\,
            I => \N__9591\
        );

    \I__2039\ : Span12Mux_v
    port map (
            O => \N__9594\,
            I => \N__9586\
        );

    \I__2038\ : Span12Mux_s10_v
    port map (
            O => \N__9591\,
            I => \N__9583\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9580\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__9589\,
            I => \N__9577\
        );

    \I__2035\ : Span12Mux_h
    port map (
            O => \N__9586\,
            I => \N__9574\
        );

    \I__2034\ : Span12Mux_h
    port map (
            O => \N__9583\,
            I => \N__9569\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9580\,
            I => \N__9569\
        );

    \I__2032\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9566\
        );

    \I__2031\ : Odrv12
    port map (
            O => \N__9574\,
            I => \TACK_EN\
        );

    \I__2030\ : Odrv12
    port map (
            O => \N__9569\,
            I => \TACK_EN\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9566\,
            I => \TACK_EN\
        );

    \I__2028\ : IoInMux
    port map (
            O => \N__9559\,
            I => \N__9556\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9556\,
            I => \N__9553\
        );

    \I__2026\ : Span4Mux_s1_v
    port map (
            O => \N__9553\,
            I => \N__9550\
        );

    \I__2025\ : Sp12to4
    port map (
            O => \N__9550\,
            I => \N__9547\
        );

    \I__2024\ : Span12Mux_s9_h
    port map (
            O => \N__9547\,
            I => \N__9544\
        );

    \I__2023\ : Span12Mux_v
    port map (
            O => \N__9544\,
            I => \N__9541\
        );

    \I__2022\ : Odrv12
    port map (
            O => \N__9541\,
            I => \TCIn_1_i\
        );

    \I__2021\ : IoInMux
    port map (
            O => \N__9538\,
            I => \N__9535\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__9535\,
            I => \N__9532\
        );

    \I__2019\ : Odrv12
    port map (
            O => \N__9532\,
            I => \RESETn_c_i\
        );

    \I__2018\ : InMux
    port map (
            O => \N__9529\,
            I => \N__9526\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__9526\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\
        );

    \I__2016\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9519\
        );

    \I__2015\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9516\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__9519\,
            I => \N__9513\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__9516\,
            I => \AC_TACK\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__9513\,
            I => \AC_TACK\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__9508\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__9505\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__9502\,
            I => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\
        );

    \I__2008\ : IoInMux
    port map (
            O => \N__9499\,
            I => \N__9495\
        );

    \I__2007\ : IoInMux
    port map (
            O => \N__9498\,
            I => \N__9492\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__9495\,
            I => \N__9486\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__9492\,
            I => \N__9486\
        );

    \I__2004\ : IoInMux
    port map (
            O => \N__9491\,
            I => \N__9483\
        );

    \I__2003\ : Span12Mux_s6_v
    port map (
            O => \N__9486\,
            I => \N__9480\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__9483\,
            I => \N__9477\
        );

    \I__2001\ : Span12Mux_v
    port map (
            O => \N__9480\,
            I => \N__9474\
        );

    \I__2000\ : Span12Mux_s11_v
    port map (
            O => \N__9477\,
            I => \N__9471\
        );

    \I__1999\ : Span12Mux_h
    port map (
            O => \N__9474\,
            I => \N__9466\
        );

    \I__1998\ : Span12Mux_h
    port map (
            O => \N__9471\,
            I => \N__9463\
        );

    \I__1997\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9458\
        );

    \I__1996\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9458\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__9466\,
            I => \TACK_OUTn\
        );

    \I__1994\ : Odrv12
    port map (
            O => \N__9463\,
            I => \TACK_OUTn\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__9458\,
            I => \TACK_OUTn\
        );

    \I__1992\ : InMux
    port map (
            O => \N__9451\,
            I => \N__9445\
        );

    \I__1991\ : InMux
    port map (
            O => \N__9450\,
            I => \N__9438\
        );

    \I__1990\ : InMux
    port map (
            O => \N__9449\,
            I => \N__9438\
        );

    \I__1989\ : InMux
    port map (
            O => \N__9448\,
            I => \N__9438\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__9445\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__9438\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\
        );

    \I__1986\ : InMux
    port map (
            O => \N__9433\,
            I => \N__9427\
        );

    \I__1985\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9420\
        );

    \I__1984\ : InMux
    port map (
            O => \N__9431\,
            I => \N__9420\
        );

    \I__1983\ : InMux
    port map (
            O => \N__9430\,
            I => \N__9420\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__9427\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__9420\,
            I => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\
        );

    \I__1980\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9411\
        );

    \I__1979\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9408\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__9411\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__9408\,
            I => \U409_TRANSFER_ACK.TACK_COUNTER6\
        );

    \I__1976\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9400\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9392\
        );

    \I__1974\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9389\
        );

    \I__1973\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9385\
        );

    \I__1972\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9382\
        );

    \I__1971\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9379\
        );

    \I__1970\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9376\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__9392\,
            I => \N__9370\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__9389\,
            I => \N__9370\
        );

    \I__1967\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9367\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__9385\,
            I => \N__9364\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9359\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__9379\,
            I => \N__9359\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__9376\,
            I => \N__9356\
        );

    \I__1962\ : InMux
    port map (
            O => \N__9375\,
            I => \N__9353\
        );

    \I__1961\ : Span4Mux_h
    port map (
            O => \N__9370\,
            I => \N__9347\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__9367\,
            I => \N__9347\
        );

    \I__1959\ : Span4Mux_v
    port map (
            O => \N__9364\,
            I => \N__9340\
        );

    \I__1958\ : Span4Mux_h
    port map (
            O => \N__9359\,
            I => \N__9340\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__9356\,
            I => \N__9340\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__9353\,
            I => \N__9337\
        );

    \I__1955\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9334\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__9347\,
            I => \N__9331\
        );

    \I__1953\ : Span4Mux_h
    port map (
            O => \N__9340\,
            I => \N__9324\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__9337\,
            I => \N__9324\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__9334\,
            I => \N__9324\
        );

    \I__1950\ : Sp12to4
    port map (
            O => \N__9331\,
            I => \N__9321\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__9324\,
            I => \N__9318\
        );

    \I__1948\ : Span12Mux_h
    port map (
            O => \N__9321\,
            I => \N__9315\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__9318\,
            I => \N__9312\
        );

    \I__1946\ : Odrv12
    port map (
            O => \N__9315\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__9312\,
            I => \U409_ADDRESS_DECODE.Z2_SPACE\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__9307\,
            I => \ROMEN_cascade_\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__9304\,
            I => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_\
        );

    \I__1942\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9293\
        );

    \I__1940\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9288\
        );

    \I__1939\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9288\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__9293\,
            I => \N__9285\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__9288\,
            I => \N__9280\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__9285\,
            I => \N__9277\
        );

    \I__1935\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9274\
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__9283\,
            I => \N__9271\
        );

    \I__1933\ : Span4Mux_h
    port map (
            O => \N__9280\,
            I => \N__9268\
        );

    \I__1932\ : Span4Mux_h
    port map (
            O => \N__9277\,
            I => \N__9263\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__9274\,
            I => \N__9263\
        );

    \I__1930\ : InMux
    port map (
            O => \N__9271\,
            I => \N__9260\
        );

    \I__1929\ : Span4Mux_h
    port map (
            O => \N__9268\,
            I => \N__9255\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__9263\,
            I => \N__9255\
        );

    \I__1927\ : LocalMux
    port map (
            O => \N__9260\,
            I => \N__9252\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__9255\,
            I => \N__9249\
        );

    \I__1925\ : Sp12to4
    port map (
            O => \N__9252\,
            I => \N__9246\
        );

    \I__1924\ : Sp12to4
    port map (
            O => \N__9249\,
            I => \N__9241\
        );

    \I__1923\ : Span12Mux_v
    port map (
            O => \N__9246\,
            I => \N__9241\
        );

    \I__1922\ : Odrv12
    port map (
            O => \N__9241\,
            I => \A_c_16\
        );

    \I__1921\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__1920\ : InMux
    port map (
            O => \N__9237\,
            I => \N__9232\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__1918\ : Span4Mux_v
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__1917\ : Sp12to4
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__1916\ : Span12Mux_h
    port map (
            O => \N__9223\,
            I => \N__9220\
        );

    \I__1915\ : Odrv12
    port map (
            O => \N__9220\,
            I => \A_c_15\
        );

    \I__1914\ : InMux
    port map (
            O => \N__9217\,
            I => \N__9212\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__9216\,
            I => \N__9209\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__9215\,
            I => \N__9206\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__9212\,
            I => \N__9203\
        );

    \I__1910\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9198\
        );

    \I__1909\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9198\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__9203\,
            I => \N__9193\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__9198\,
            I => \N__9193\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__1905\ : Sp12to4
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__1904\ : Span12Mux_h
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__1903\ : Odrv12
    port map (
            O => \N__9184\,
            I => \A_c_13\
        );

    \I__1902\ : IoInMux
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__9178\,
            I => \N__9175\
        );

    \I__1900\ : IoSpan4Mux
    port map (
            O => \N__9175\,
            I => \N__9172\
        );

    \I__1899\ : Span4Mux_s2_h
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__1898\ : Sp12to4
    port map (
            O => \N__9169\,
            I => \N__9166\
        );

    \I__1897\ : Span12Mux_h
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__1896\ : Odrv12
    port map (
            O => \N__9163\,
            I => \U409_ADDRESS_DECODE_un1_CIACS1n_i\
        );

    \I__1895\ : InMux
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__9157\,
            I => \CIA_ENABLE\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \CIA_ENABLE_cascade_\
        );

    \I__1892\ : InMux
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__1891\ : InMux
    port map (
            O => \N__9150\,
            I => \N__9145\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__9145\,
            I => \N__9142\
        );

    \I__1889\ : Span4Mux_v
    port map (
            O => \N__9142\,
            I => \N__9138\
        );

    \I__1888\ : InMux
    port map (
            O => \N__9141\,
            I => \N__9135\
        );

    \I__1887\ : Sp12to4
    port map (
            O => \N__9138\,
            I => \N__9130\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__9135\,
            I => \N__9130\
        );

    \I__1885\ : Span12Mux_h
    port map (
            O => \N__9130\,
            I => \N__9127\
        );

    \I__1884\ : Odrv12
    port map (
            O => \N__9127\,
            I => \A_c_12\
        );

    \I__1883\ : IoInMux
    port map (
            O => \N__9124\,
            I => \N__9121\
        );

    \I__1882\ : LocalMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__1881\ : IoSpan4Mux
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__1880\ : IoSpan4Mux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__1879\ : Span4Mux_s3_h
    port map (
            O => \N__9112\,
            I => \N__9109\
        );

    \I__1878\ : Span4Mux_h
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__1877\ : Sp12to4
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__1876\ : Odrv12
    port map (
            O => \N__9103\,
            I => \U409_ADDRESS_DECODE_un1_CIACS0n_i\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__1874\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9093\
        );

    \I__1873\ : InMux
    port map (
            O => \N__9096\,
            I => \N__9089\
        );

    \I__1872\ : LocalMux
    port map (
            O => \N__9093\,
            I => \N__9086\
        );

    \I__1871\ : InMux
    port map (
            O => \N__9092\,
            I => \N__9083\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__9089\,
            I => \N__9079\
        );

    \I__1869\ : Span4Mux_v
    port map (
            O => \N__9086\,
            I => \N__9076\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__9083\,
            I => \N__9073\
        );

    \I__1867\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9070\
        );

    \I__1866\ : Span12Mux_v
    port map (
            O => \N__9079\,
            I => \N__9067\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__9076\,
            I => \N__9064\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__9073\,
            I => \N__9061\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__9070\,
            I => \N__9058\
        );

    \I__1862\ : Odrv12
    port map (
            O => \N__9067\,
            I => \U409_ADDRESS_DECODE.N_75\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__9064\,
            I => \U409_ADDRESS_DECODE.N_75\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__9061\,
            I => \U409_ADDRESS_DECODE.N_75\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__9058\,
            I => \U409_ADDRESS_DECODE.N_75\
        );

    \I__1858\ : IoInMux
    port map (
            O => \N__9049\,
            I => \N__9046\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__1856\ : Span4Mux_s3_h
    port map (
            O => \N__9043\,
            I => \N__9040\
        );

    \I__1855\ : Span4Mux_v
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__1854\ : Span4Mux_h
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__1853\ : Span4Mux_h
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__1852\ : Span4Mux_h
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__1851\ : Odrv4
    port map (
            O => \N__9028\,
            I => \N_77_mux_i\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \N__9022\
        );

    \I__1849\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9019\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__9019\,
            I => \N__9015\
        );

    \I__1847\ : InMux
    port map (
            O => \N__9018\,
            I => \N__9012\
        );

    \I__1846\ : Span4Mux_v
    port map (
            O => \N__9015\,
            I => \N__9009\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__9012\,
            I => \N__9006\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__9009\,
            I => \U409_ADDRESS_DECODE.N_60_1\
        );

    \I__1843\ : Odrv4
    port map (
            O => \N__9006\,
            I => \U409_ADDRESS_DECODE.N_60_1\
        );

    \I__1842\ : IoInMux
    port map (
            O => \N__9001\,
            I => \N__8998\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__1840\ : Span12Mux_s11_v
    port map (
            O => \N__8995\,
            I => \N__8992\
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__8992\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\
        );

    \I__1838\ : InMux
    port map (
            O => \N__8989\,
            I => \N__8986\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__1836\ : Odrv4
    port map (
            O => \N__8983\,
            I => \U409_AUTOCONFIG.STATE4\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8973\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8968\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8968\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8965\
        );

    \I__1831\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8962\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__8973\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__8968\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8965\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8962\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__8953\,
            I => \N__8950\
        );

    \I__1825\ : InMux
    port map (
            O => \N__8950\,
            I => \N__8947\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8947\,
            I => \N_71_mux\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8939\
        );

    \I__1822\ : InMux
    port map (
            O => \N__8943\,
            I => \N__8936\
        );

    \I__1821\ : InMux
    port map (
            O => \N__8942\,
            I => \N__8933\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8939\,
            I => \N_70_mux\
        );

    \I__1819\ : LocalMux
    port map (
            O => \N__8936\,
            I => \N_70_mux\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__8933\,
            I => \N_70_mux\
        );

    \I__1817\ : CEMux
    port map (
            O => \N__8926\,
            I => \N__8923\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__8923\,
            I => \U409_TRANSFER_ACK.N_20_0\
        );

    \I__1815\ : InMux
    port map (
            O => \N__8920\,
            I => \N__8916\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8913\
        );

    \I__1813\ : LocalMux
    port map (
            O => \N__8916\,
            I => \N__8910\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__8913\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__8910\,
            I => \U409_AUTOCONFIG.STATE_d_2\
        );

    \I__1810\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1809\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8896\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__8903\,
            I => \N__8892\
        );

    \I__1807\ : InMux
    port map (
            O => \N__8902\,
            I => \N__8888\
        );

    \I__1806\ : LocalMux
    port map (
            O => \N__8899\,
            I => \N__8883\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__8896\,
            I => \N__8883\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8876\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8892\,
            I => \N__8876\
        );

    \I__1802\ : InMux
    port map (
            O => \N__8891\,
            I => \N__8876\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8888\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1800\ : Odrv12
    port map (
            O => \N__8883\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__8876\,
            I => \U409_AUTOCONFIG.STATEZ0Z_1\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8868\,
            I => \N__8860\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8867\,
            I => \N__8857\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8866\,
            I => \N__8853\
        );

    \I__1794\ : InMux
    port map (
            O => \N__8863\,
            I => \N__8850\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8860\,
            I => \N__8847\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8857\,
            I => \N__8844\
        );

    \I__1791\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8841\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8853\,
            I => \N__8838\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__8850\,
            I => \N__8834\
        );

    \I__1788\ : Span4Mux_v
    port map (
            O => \N__8847\,
            I => \N__8831\
        );

    \I__1787\ : Span4Mux_v
    port map (
            O => \N__8844\,
            I => \N__8826\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__8841\,
            I => \N__8826\
        );

    \I__1785\ : Span4Mux_v
    port map (
            O => \N__8838\,
            I => \N__8823\
        );

    \I__1784\ : InMux
    port map (
            O => \N__8837\,
            I => \N__8820\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__8834\,
            I => \N__8817\
        );

    \I__1782\ : Span4Mux_v
    port map (
            O => \N__8831\,
            I => \N__8814\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__8826\,
            I => \N__8811\
        );

    \I__1780\ : Sp12to4
    port map (
            O => \N__8823\,
            I => \N__8806\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__8820\,
            I => \N__8806\
        );

    \I__1778\ : Sp12to4
    port map (
            O => \N__8817\,
            I => \N__8799\
        );

    \I__1777\ : Sp12to4
    port map (
            O => \N__8814\,
            I => \N__8799\
        );

    \I__1776\ : Sp12to4
    port map (
            O => \N__8811\,
            I => \N__8799\
        );

    \I__1775\ : Span12Mux_h
    port map (
            O => \N__8806\,
            I => \N__8796\
        );

    \I__1774\ : Span12Mux_h
    port map (
            O => \N__8799\,
            I => \N__8793\
        );

    \I__1773\ : Span12Mux_v
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__1772\ : Span12Mux_v
    port map (
            O => \N__8793\,
            I => \N__8787\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__8790\,
            I => \RnW_c\
        );

    \I__1770\ : Odrv12
    port map (
            O => \N__8787\,
            I => \RnW_c\
        );

    \I__1769\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8779\
        );

    \I__1768\ : LocalMux
    port map (
            O => \N__8779\,
            I => \N__8774\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8771\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8765\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__8774\,
            I => \N__8762\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8771\,
            I => \N__8759\
        );

    \I__1763\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8752\
        );

    \I__1762\ : InMux
    port map (
            O => \N__8769\,
            I => \N__8752\
        );

    \I__1761\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8752\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__8765\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1759\ : Odrv4
    port map (
            O => \N__8762\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1758\ : Odrv12
    port map (
            O => \N__8759\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__8752\,
            I => \U409_AUTOCONFIG.STATEZ0Z_0\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8743\,
            I => \N__8739\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8742\,
            I => \N__8736\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8733\
        );

    \I__1753\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8730\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8733\,
            I => \N__8727\
        );

    \I__1751\ : Span4Mux_v
    port map (
            O => \N__8730\,
            I => \N__8723\
        );

    \I__1750\ : Span4Mux_v
    port map (
            O => \N__8727\,
            I => \N__8720\
        );

    \I__1749\ : InMux
    port map (
            O => \N__8726\,
            I => \N__8717\
        );

    \I__1748\ : Odrv4
    port map (
            O => \N__8723\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1747\ : Odrv4
    port map (
            O => \N__8720\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__8717\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8707\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__8707\,
            I => \N__8704\
        );

    \I__1743\ : Sp12to4
    port map (
            O => \N__8704\,
            I => \N__8701\
        );

    \I__1742\ : Span12Mux_v
    port map (
            O => \N__8701\,
            I => \N__8698\
        );

    \I__1741\ : Span12Mux_h
    port map (
            O => \N__8698\,
            I => \N__8695\
        );

    \I__1740\ : Odrv12
    port map (
            O => \N__8695\,
            I => \TACKn_in\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__8692\,
            I => \N__8689\
        );

    \I__1738\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8685\
        );

    \I__1737\ : InMux
    port map (
            O => \N__8688\,
            I => \N__8682\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__8685\,
            I => \N__8677\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__8682\,
            I => \N__8677\
        );

    \I__1734\ : Odrv12
    port map (
            O => \N__8677\,
            I => \U409_ADDRESS_DECODE_un1_RAMSPACEn\
        );

    \I__1733\ : SRMux
    port map (
            O => \N__8674\,
            I => \N__8670\
        );

    \I__1732\ : SRMux
    port map (
            O => \N__8673\,
            I => \N__8667\
        );

    \I__1731\ : LocalMux
    port map (
            O => \N__8670\,
            I => \N__8663\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8667\,
            I => \N__8660\
        );

    \I__1729\ : SRMux
    port map (
            O => \N__8666\,
            I => \N__8657\
        );

    \I__1728\ : Span4Mux_v
    port map (
            O => \N__8663\,
            I => \N__8651\
        );

    \I__1727\ : Span4Mux_h
    port map (
            O => \N__8660\,
            I => \N__8651\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__8657\,
            I => \N__8648\
        );

    \I__1725\ : SRMux
    port map (
            O => \N__8656\,
            I => \N__8645\
        );

    \I__1724\ : Odrv4
    port map (
            O => \N__8651\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__8648\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__8645\,
            I => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\
        );

    \I__1721\ : IoInMux
    port map (
            O => \N__8638\,
            I => \N__8635\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8632\
        );

    \I__1719\ : Span4Mux_s2_v
    port map (
            O => \N__8632\,
            I => \N__8629\
        );

    \I__1718\ : Span4Mux_v
    port map (
            O => \N__8629\,
            I => \N__8626\
        );

    \I__1717\ : Odrv4
    port map (
            O => \N__8626\,
            I => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__8623\,
            I => \N__8616\
        );

    \I__1715\ : InMux
    port map (
            O => \N__8622\,
            I => \N__8609\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8609\
        );

    \I__1713\ : InMux
    port map (
            O => \N__8620\,
            I => \N__8609\
        );

    \I__1712\ : InMux
    port map (
            O => \N__8619\,
            I => \N__8604\
        );

    \I__1711\ : InMux
    port map (
            O => \N__8616\,
            I => \N__8604\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N_23\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N_23\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__8599\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__8596\,
            I => \N__8592\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__8595\,
            I => \N__8587\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8592\,
            I => \N__8579\
        );

    \I__1704\ : InMux
    port map (
            O => \N__8591\,
            I => \N__8579\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8590\,
            I => \N__8579\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8587\,
            I => \N__8574\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8586\,
            I => \N__8574\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__8579\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__8574\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3\
        );

    \I__1698\ : InMux
    port map (
            O => \N__8569\,
            I => \N__8560\
        );

    \I__1697\ : InMux
    port map (
            O => \N__8568\,
            I => \N__8560\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8567\,
            I => \N__8553\
        );

    \I__1695\ : InMux
    port map (
            O => \N__8566\,
            I => \N__8553\
        );

    \I__1694\ : InMux
    port map (
            O => \N__8565\,
            I => \N__8553\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__8560\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8553\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8545\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8545\,
            I => \N__8539\
        );

    \I__1689\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8536\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8533\
        );

    \I__1687\ : InMux
    port map (
            O => \N__8542\,
            I => \N__8529\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__8539\,
            I => \N__8524\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__8536\,
            I => \N__8524\
        );

    \I__1684\ : LocalMux
    port map (
            O => \N__8533\,
            I => \N__8521\
        );

    \I__1683\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8518\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8515\
        );

    \I__1681\ : Span4Mux_v
    port map (
            O => \N__8524\,
            I => \N__8508\
        );

    \I__1680\ : Span4Mux_v
    port map (
            O => \N__8521\,
            I => \N__8508\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__8518\,
            I => \N__8508\
        );

    \I__1678\ : Odrv12
    port map (
            O => \N__8515\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_4\
        );

    \I__1677\ : Odrv4
    port map (
            O => \N__8508\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_4\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__8503\,
            I => \N__8500\
        );

    \I__1675\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8497\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8492\
        );

    \I__1673\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8489\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__8495\,
            I => \N__8486\
        );

    \I__1671\ : Span4Mux_v
    port map (
            O => \N__8492\,
            I => \N__8481\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__8489\,
            I => \N__8481\
        );

    \I__1669\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8478\
        );

    \I__1668\ : Span4Mux_h
    port map (
            O => \N__8481\,
            I => \N__8474\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__8478\,
            I => \N__8471\
        );

    \I__1666\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8468\
        );

    \I__1665\ : Span4Mux_v
    port map (
            O => \N__8474\,
            I => \N__8463\
        );

    \I__1664\ : Span4Mux_v
    port map (
            O => \N__8471\,
            I => \N__8463\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__8468\,
            I => \N__8460\
        );

    \I__1662\ : Odrv4
    port map (
            O => \N__8463\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_5\
        );

    \I__1661\ : Odrv12
    port map (
            O => \N__8460\,
            I => \U409_ADDRESS_DECODE.CIA_SPACE_5\
        );

    \I__1660\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8451\
        );

    \I__1659\ : InMux
    port map (
            O => \N__8454\,
            I => \N__8448\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__8451\,
            I => \LIDE_BASE_4\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__8448\,
            I => \LIDE_BASE_4\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__8443\,
            I => \N__8440\
        );

    \I__1655\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8436\
        );

    \I__1654\ : InMux
    port map (
            O => \N__8439\,
            I => \N__8433\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__8436\,
            I => \LIDE_BASE_3\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__8433\,
            I => \LIDE_BASE_3\
        );

    \I__1651\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8425\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__8425\,
            I => \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\
        );

    \I__1649\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8418\
        );

    \I__1648\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8414\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8410\
        );

    \I__1646\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8407\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8404\
        );

    \I__1644\ : InMux
    port map (
            O => \N__8413\,
            I => \N__8401\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__8410\,
            I => \N__8398\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__8407\,
            I => \N__8391\
        );

    \I__1641\ : Span4Mux_v
    port map (
            O => \N__8404\,
            I => \N__8391\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__8401\,
            I => \N__8391\
        );

    \I__1639\ : Span4Mux_h
    port map (
            O => \N__8398\,
            I => \N__8385\
        );

    \I__1638\ : Span4Mux_v
    port map (
            O => \N__8391\,
            I => \N__8385\
        );

    \I__1637\ : InMux
    port map (
            O => \N__8390\,
            I => \N__8382\
        );

    \I__1636\ : Odrv4
    port map (
            O => \N__8385\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__8382\,
            I => \AUTOCONFIG_SPACE\
        );

    \I__1634\ : IoInMux
    port map (
            O => \N__8377\,
            I => \N__8374\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__8374\,
            I => \N__8371\
        );

    \I__1632\ : Span12Mux_s7_v
    port map (
            O => \N__8371\,
            I => \N__8368\
        );

    \I__1631\ : Span12Mux_v
    port map (
            O => \N__8368\,
            I => \N__8365\
        );

    \I__1630\ : Odrv12
    port map (
            O => \N__8365\,
            I => \BUFENn_c\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__8362\,
            I => \N__8359\
        );

    \I__1628\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8352\
        );

    \I__1627\ : InMux
    port map (
            O => \N__8358\,
            I => \N__8352\
        );

    \I__1626\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8349\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__8352\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__8349\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0\
        );

    \I__1623\ : InMux
    port map (
            O => \N__8344\,
            I => \N__8339\
        );

    \I__1622\ : InMux
    port map (
            O => \N__8343\,
            I => \N__8334\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8334\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__8339\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8334\,
            I => \U409_ADDRESS_DECODE.ATA_ENZ0\
        );

    \I__1618\ : IoInMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8323\
        );

    \I__1616\ : IoSpan4Mux
    port map (
            O => \N__8323\,
            I => \N__8320\
        );

    \I__1615\ : Sp12to4
    port map (
            O => \N__8320\,
            I => \N__8317\
        );

    \I__1614\ : Span12Mux_s7_h
    port map (
            O => \N__8317\,
            I => \N__8314\
        );

    \I__1613\ : Odrv12
    port map (
            O => \N__8314\,
            I => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__1611\ : InMux
    port map (
            O => \N__8310\,
            I => \N__8302\
        );

    \I__1610\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8299\
        );

    \I__1609\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8294\
        );

    \I__1608\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8294\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__8302\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__8299\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__8294\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__8287\,
            I => \U409_ADDRESS_DECODE.m27Z0Z_3_cascade_\
        );

    \I__1603\ : InMux
    port map (
            O => \N__8284\,
            I => \N__8278\
        );

    \I__1602\ : InMux
    port map (
            O => \N__8283\,
            I => \N__8278\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__8278\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__8275\,
            I => \N__8270\
        );

    \I__1599\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8264\
        );

    \I__1598\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8264\
        );

    \I__1597\ : InMux
    port map (
            O => \N__8270\,
            I => \N__8259\
        );

    \I__1596\ : InMux
    port map (
            O => \N__8269\,
            I => \N__8259\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__8264\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__8259\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4\
        );

    \I__1593\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8251\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__8251\,
            I => \U409_ADDRESS_DECODE_m33_1\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__8248\,
            I => \U409_ADDRESS_DECODE_m33_1_cascade_\
        );

    \I__1590\ : InMux
    port map (
            O => \N__8245\,
            I => \N__8239\
        );

    \I__1589\ : InMux
    port map (
            O => \N__8244\,
            I => \N__8236\
        );

    \I__1588\ : InMux
    port map (
            O => \N__8243\,
            I => \N__8231\
        );

    \I__1587\ : InMux
    port map (
            O => \N__8242\,
            I => \N__8231\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__8239\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5\
        );

    \I__1585\ : LocalMux
    port map (
            O => \N__8236\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__8231\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5\
        );

    \I__1583\ : InMux
    port map (
            O => \N__8224\,
            I => \N__8218\
        );

    \I__1582\ : InMux
    port map (
            O => \N__8223\,
            I => \N__8211\
        );

    \I__1581\ : InMux
    port map (
            O => \N__8222\,
            I => \N__8211\
        );

    \I__1580\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8211\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__8218\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__8211\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__8206\,
            I => \N__8202\
        );

    \I__1576\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8199\
        );

    \I__1575\ : InMux
    port map (
            O => \N__8202\,
            I => \N__8196\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__8199\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__8196\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2\
        );

    \I__1572\ : InMux
    port map (
            O => \N__8191\,
            I => \N__8184\
        );

    \I__1571\ : InMux
    port map (
            O => \N__8190\,
            I => \N__8181\
        );

    \I__1570\ : InMux
    port map (
            O => \N__8189\,
            I => \N__8178\
        );

    \I__1569\ : InMux
    port map (
            O => \N__8188\,
            I => \N__8173\
        );

    \I__1568\ : InMux
    port map (
            O => \N__8187\,
            I => \N__8173\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__8184\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__8181\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__8178\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__8173\,
            I => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__8164\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_\
        );

    \I__1562\ : InMux
    port map (
            O => \N__8161\,
            I => \N__8155\
        );

    \I__1561\ : InMux
    port map (
            O => \N__8160\,
            I => \N__8155\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__8155\,
            I => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__8152\,
            I => \N__8149\
        );

    \I__1558\ : InMux
    port map (
            O => \N__8149\,
            I => \N__8144\
        );

    \I__1557\ : InMux
    port map (
            O => \N__8148\,
            I => \N__8139\
        );

    \I__1556\ : InMux
    port map (
            O => \N__8147\,
            I => \N__8139\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__8144\,
            I => \N__8134\
        );

    \I__1554\ : LocalMux
    port map (
            O => \N__8139\,
            I => \N__8131\
        );

    \I__1553\ : CascadeMux
    port map (
            O => \N__8138\,
            I => \N__8128\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__8137\,
            I => \N__8125\
        );

    \I__1551\ : Span4Mux_v
    port map (
            O => \N__8134\,
            I => \N__8120\
        );

    \I__1550\ : Span4Mux_v
    port map (
            O => \N__8131\,
            I => \N__8120\
        );

    \I__1549\ : InMux
    port map (
            O => \N__8128\,
            I => \N__8115\
        );

    \I__1548\ : InMux
    port map (
            O => \N__8125\,
            I => \N__8115\
        );

    \I__1547\ : Sp12to4
    port map (
            O => \N__8120\,
            I => \N__8110\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8110\
        );

    \I__1545\ : Span12Mux_h
    port map (
            O => \N__8110\,
            I => \N__8107\
        );

    \I__1544\ : Span12Mux_v
    port map (
            O => \N__8107\,
            I => \N__8104\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__8104\,
            I => \D_in_5\
        );

    \I__1542\ : InMux
    port map (
            O => \N__8101\,
            I => \N__8098\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__8098\,
            I => \N__8094\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__8097\,
            I => \N__8091\
        );

    \I__1539\ : Span4Mux_v
    port map (
            O => \N__8094\,
            I => \N__8088\
        );

    \I__1538\ : InMux
    port map (
            O => \N__8091\,
            I => \N__8085\
        );

    \I__1537\ : Odrv4
    port map (
            O => \N__8088\,
            I => \BRIDGE_BASE_1\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__8085\,
            I => \BRIDGE_BASE_1\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__8080\,
            I => \N__8077\
        );

    \I__1534\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8073\
        );

    \I__1533\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8070\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__8073\,
            I => \N__8067\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__8070\,
            I => \LIDE_BASE_7\
        );

    \I__1530\ : Odrv12
    port map (
            O => \N__8067\,
            I => \LIDE_BASE_7\
        );

    \I__1529\ : CascadeMux
    port map (
            O => \N__8062\,
            I => \N__8058\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__8061\,
            I => \N__8055\
        );

    \I__1527\ : InMux
    port map (
            O => \N__8058\,
            I => \N__8052\
        );

    \I__1526\ : InMux
    port map (
            O => \N__8055\,
            I => \N__8049\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__8052\,
            I => \N__8043\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__8049\,
            I => \N__8040\
        );

    \I__1523\ : InMux
    port map (
            O => \N__8048\,
            I => \N__8033\
        );

    \I__1522\ : InMux
    port map (
            O => \N__8047\,
            I => \N__8033\
        );

    \I__1521\ : InMux
    port map (
            O => \N__8046\,
            I => \N__8033\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__8043\,
            I => \N__8030\
        );

    \I__1519\ : Span4Mux_h
    port map (
            O => \N__8040\,
            I => \N__8025\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__8033\,
            I => \N__8025\
        );

    \I__1517\ : Span4Mux_h
    port map (
            O => \N__8030\,
            I => \N__8020\
        );

    \I__1516\ : Span4Mux_v
    port map (
            O => \N__8025\,
            I => \N__8020\
        );

    \I__1515\ : Sp12to4
    port map (
            O => \N__8020\,
            I => \N__8017\
        );

    \I__1514\ : Odrv12
    port map (
            O => \N__8017\,
            I => \D_in_7\
        );

    \I__1513\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8008\
        );

    \I__1512\ : InMux
    port map (
            O => \N__8013\,
            I => \N__8003\
        );

    \I__1511\ : InMux
    port map (
            O => \N__8012\,
            I => \N__8003\
        );

    \I__1510\ : InMux
    port map (
            O => \N__8011\,
            I => \N__8000\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__8008\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__8003\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__8000\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__7993\,
            I => \N__7990\
        );

    \I__1505\ : InMux
    port map (
            O => \N__7990\,
            I => \N__7986\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__7989\,
            I => \N__7983\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__7986\,
            I => \N__7980\
        );

    \I__1502\ : InMux
    port map (
            O => \N__7983\,
            I => \N__7977\
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__7980\,
            I => \BRIDGE_BASE_3\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7977\,
            I => \BRIDGE_BASE_3\
        );

    \I__1499\ : InMux
    port map (
            O => \N__7972\,
            I => \N__7964\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7971\,
            I => \N__7964\
        );

    \I__1497\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7959\
        );

    \I__1496\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7959\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__7964\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7959\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__7954\,
            I => \N__7949\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__7953\,
            I => \N__7946\
        );

    \I__1491\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7943\
        );

    \I__1490\ : InMux
    port map (
            O => \N__7949\,
            I => \N__7940\
        );

    \I__1489\ : InMux
    port map (
            O => \N__7946\,
            I => \N__7937\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__7943\,
            I => \N__7930\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__7940\,
            I => \N__7930\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__7937\,
            I => \N__7930\
        );

    \I__1485\ : Span4Mux_v
    port map (
            O => \N__7930\,
            I => \N__7927\
        );

    \I__1484\ : Sp12to4
    port map (
            O => \N__7927\,
            I => \N__7924\
        );

    \I__1483\ : Span12Mux_h
    port map (
            O => \N__7924\,
            I => \N__7921\
        );

    \I__1482\ : Odrv12
    port map (
            O => \N__7921\,
            I => \D_in_4\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7918\,
            I => \N__7914\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__7917\,
            I => \N__7911\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7914\,
            I => \N__7891\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7911\,
            I => \N__7891\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7891\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7891\
        );

    \I__1475\ : InMux
    port map (
            O => \N__7908\,
            I => \N__7891\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7907\,
            I => \N__7891\
        );

    \I__1473\ : InMux
    port map (
            O => \N__7906\,
            I => \N__7881\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7881\
        );

    \I__1471\ : InMux
    port map (
            O => \N__7904\,
            I => \N__7881\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7891\,
            I => \N__7878\
        );

    \I__1469\ : InMux
    port map (
            O => \N__7890\,
            I => \N__7866\
        );

    \I__1468\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7866\
        );

    \I__1467\ : InMux
    port map (
            O => \N__7888\,
            I => \N__7866\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7881\,
            I => \N__7862\
        );

    \I__1465\ : Span4Mux_v
    port map (
            O => \N__7878\,
            I => \N__7859\
        );

    \I__1464\ : InMux
    port map (
            O => \N__7877\,
            I => \N__7854\
        );

    \I__1463\ : InMux
    port map (
            O => \N__7876\,
            I => \N__7854\
        );

    \I__1462\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7847\
        );

    \I__1461\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7847\
        );

    \I__1460\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7847\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__7866\,
            I => \N__7844\
        );

    \I__1458\ : InMux
    port map (
            O => \N__7865\,
            I => \N__7841\
        );

    \I__1457\ : Span4Mux_v
    port map (
            O => \N__7862\,
            I => \N__7832\
        );

    \I__1456\ : Span4Mux_h
    port map (
            O => \N__7859\,
            I => \N__7832\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__7854\,
            I => \N__7832\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__7847\,
            I => \N__7832\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__7844\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__7841\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__7832\,
            I => \un1_AUTOCONFIG_SPACE\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__7825\,
            I => \N_71_mux_cascade_\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__7822\,
            I => \N_23_cascade_\
        );

    \I__1448\ : InMux
    port map (
            O => \N__7819\,
            I => \N__7816\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7816\,
            I => \U409_ADDRESS_DECODE.m33Z0Z_3\
        );

    \I__1446\ : InMux
    port map (
            O => \N__7813\,
            I => \N__7810\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__7810\,
            I => \N__7806\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7809\,
            I => \N__7802\
        );

    \I__1443\ : Span4Mux_v
    port map (
            O => \N__7806\,
            I => \N__7799\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7805\,
            I => \N__7794\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7802\,
            I => \N__7791\
        );

    \I__1440\ : Sp12to4
    port map (
            O => \N__7799\,
            I => \N__7788\
        );

    \I__1439\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7783\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7783\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7780\
        );

    \I__1436\ : Span4Mux_v
    port map (
            O => \N__7791\,
            I => \N__7777\
        );

    \I__1435\ : Span12Mux_h
    port map (
            O => \N__7788\,
            I => \N__7774\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7783\,
            I => \N__7771\
        );

    \I__1433\ : Sp12to4
    port map (
            O => \N__7780\,
            I => \N__7768\
        );

    \I__1432\ : Span4Mux_v
    port map (
            O => \N__7777\,
            I => \N__7765\
        );

    \I__1431\ : Span12Mux_v
    port map (
            O => \N__7774\,
            I => \N__7762\
        );

    \I__1430\ : Span12Mux_v
    port map (
            O => \N__7771\,
            I => \N__7759\
        );

    \I__1429\ : Span12Mux_v
    port map (
            O => \N__7768\,
            I => \N__7754\
        );

    \I__1428\ : Sp12to4
    port map (
            O => \N__7765\,
            I => \N__7754\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__7762\,
            I => \A_c_18\
        );

    \I__1426\ : Odrv12
    port map (
            O => \N__7759\,
            I => \A_c_18\
        );

    \I__1425\ : Odrv12
    port map (
            O => \N__7754\,
            I => \A_c_18\
        );

    \I__1424\ : InMux
    port map (
            O => \N__7747\,
            I => \N__7743\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7746\,
            I => \N__7740\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7743\,
            I => \LIDE_BASE_1\
        );

    \I__1421\ : LocalMux
    port map (
            O => \N__7740\,
            I => \LIDE_BASE_1\
        );

    \I__1420\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7729\
        );

    \I__1419\ : InMux
    port map (
            O => \N__7734\,
            I => \N__7724\
        );

    \I__1418\ : InMux
    port map (
            O => \N__7733\,
            I => \N__7724\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7732\,
            I => \N__7720\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__7729\,
            I => \N__7717\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__7724\,
            I => \N__7714\
        );

    \I__1414\ : InMux
    port map (
            O => \N__7723\,
            I => \N__7711\
        );

    \I__1413\ : InMux
    port map (
            O => \N__7720\,
            I => \N__7707\
        );

    \I__1412\ : Span4Mux_v
    port map (
            O => \N__7717\,
            I => \N__7704\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__7714\,
            I => \N__7701\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7698\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7710\,
            I => \N__7695\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__7707\,
            I => \N__7692\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__7704\,
            I => \N__7689\
        );

    \I__1406\ : Sp12to4
    port map (
            O => \N__7701\,
            I => \N__7686\
        );

    \I__1405\ : Span4Mux_h
    port map (
            O => \N__7698\,
            I => \N__7681\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7695\,
            I => \N__7681\
        );

    \I__1403\ : Span12Mux_v
    port map (
            O => \N__7692\,
            I => \N__7678\
        );

    \I__1402\ : Span4Mux_v
    port map (
            O => \N__7689\,
            I => \N__7675\
        );

    \I__1401\ : Span12Mux_h
    port map (
            O => \N__7686\,
            I => \N__7670\
        );

    \I__1400\ : Sp12to4
    port map (
            O => \N__7681\,
            I => \N__7670\
        );

    \I__1399\ : Span12Mux_h
    port map (
            O => \N__7678\,
            I => \N__7667\
        );

    \I__1398\ : Sp12to4
    port map (
            O => \N__7675\,
            I => \N__7662\
        );

    \I__1397\ : Span12Mux_v
    port map (
            O => \N__7670\,
            I => \N__7662\
        );

    \I__1396\ : Odrv12
    port map (
            O => \N__7667\,
            I => \A_c_17\
        );

    \I__1395\ : Odrv12
    port map (
            O => \N__7662\,
            I => \A_c_17\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__7657\,
            I => \N__7654\
        );

    \I__1393\ : InMux
    port map (
            O => \N__7654\,
            I => \N__7650\
        );

    \I__1392\ : InMux
    port map (
            O => \N__7653\,
            I => \N__7647\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__7650\,
            I => \LIDE_BASE_2\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7647\,
            I => \LIDE_BASE_2\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7642\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_\
        );

    \I__1388\ : CascadeMux
    port map (
            O => \N__7639\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__7636\,
            I => \N__7632\
        );

    \I__1386\ : InMux
    port map (
            O => \N__7635\,
            I => \N__7626\
        );

    \I__1385\ : InMux
    port map (
            O => \N__7632\,
            I => \N__7626\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7631\,
            I => \N__7621\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__7626\,
            I => \N__7617\
        );

    \I__1382\ : InMux
    port map (
            O => \N__7625\,
            I => \N__7614\
        );

    \I__1381\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7609\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7605\
        );

    \I__1379\ : InMux
    port map (
            O => \N__7620\,
            I => \N__7602\
        );

    \I__1378\ : Span4Mux_h
    port map (
            O => \N__7617\,
            I => \N__7597\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__7614\,
            I => \N__7597\
        );

    \I__1376\ : InMux
    port map (
            O => \N__7613\,
            I => \N__7594\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7612\,
            I => \N__7591\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7609\,
            I => \N__7588\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7608\,
            I => \N__7585\
        );

    \I__1372\ : Odrv12
    port map (
            O => \N__7605\,
            I => \CONFIGURED\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7602\,
            I => \CONFIGURED\
        );

    \I__1370\ : Odrv4
    port map (
            O => \N__7597\,
            I => \CONFIGURED\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7594\,
            I => \CONFIGURED\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__7591\,
            I => \CONFIGURED\
        );

    \I__1367\ : Odrv4
    port map (
            O => \N__7588\,
            I => \CONFIGURED\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__7585\,
            I => \CONFIGURED\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7570\,
            I => \N__7567\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7567\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__7564\,
            I => \N__7561\
        );

    \I__1362\ : InMux
    port map (
            O => \N__7561\,
            I => \N__7557\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7560\,
            I => \N__7554\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7557\,
            I => \LIDE_BASE_6\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__7554\,
            I => \LIDE_BASE_6\
        );

    \I__1358\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7545\
        );

    \I__1357\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7542\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__7545\,
            I => \LIDE_BASE_5\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__7542\,
            I => \LIDE_BASE_5\
        );

    \I__1354\ : InMux
    port map (
            O => \N__7537\,
            I => \N__7534\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__7534\,
            I => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\
        );

    \I__1352\ : InMux
    port map (
            O => \N__7531\,
            I => \N__7526\
        );

    \I__1351\ : InMux
    port map (
            O => \N__7530\,
            I => \N__7521\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7529\,
            I => \N__7521\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__7526\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__7521\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0\
        );

    \I__1347\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7513\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7509\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7512\,
            I => \N__7506\
        );

    \I__1344\ : Span4Mux_v
    port map (
            O => \N__7509\,
            I => \N__7503\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7506\,
            I => \N__7500\
        );

    \I__1342\ : Odrv4
    port map (
            O => \N__7503\,
            I => \BRIDGE_BASE_5\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7500\,
            I => \BRIDGE_BASE_5\
        );

    \I__1340\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7490\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7494\,
            I => \N__7485\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7493\,
            I => \N__7485\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7482\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__7485\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0\
        );

    \I__1335\ : Odrv4
    port map (
            O => \N__7482\,
            I => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0\
        );

    \I__1334\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7474\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__7474\,
            I => \N__7471\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__7471\,
            I => \N__7468\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__7468\,
            I => \N__7464\
        );

    \I__1330\ : InMux
    port map (
            O => \N__7467\,
            I => \N__7461\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__7464\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_13\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__7461\,
            I => \U409_AUTOCONFIG.un1_AZ0Z_13\
        );

    \I__1327\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7452\
        );

    \I__1326\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7445\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__7452\,
            I => \N__7442\
        );

    \I__1324\ : InMux
    port map (
            O => \N__7451\,
            I => \N__7439\
        );

    \I__1323\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7432\
        );

    \I__1322\ : InMux
    port map (
            O => \N__7449\,
            I => \N__7429\
        );

    \I__1321\ : InMux
    port map (
            O => \N__7448\,
            I => \N__7424\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7417\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__7442\,
            I => \N__7417\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__7439\,
            I => \N__7417\
        );

    \I__1317\ : InMux
    port map (
            O => \N__7438\,
            I => \N__7408\
        );

    \I__1316\ : InMux
    port map (
            O => \N__7437\,
            I => \N__7408\
        );

    \I__1315\ : InMux
    port map (
            O => \N__7436\,
            I => \N__7408\
        );

    \I__1314\ : InMux
    port map (
            O => \N__7435\,
            I => \N__7408\
        );

    \I__1313\ : InMux
    port map (
            O => \N__7432\,
            I => \N__7403\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7400\
        );

    \I__1311\ : InMux
    port map (
            O => \N__7428\,
            I => \N__7397\
        );

    \I__1310\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7394\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__7424\,
            I => \N__7387\
        );

    \I__1308\ : Span4Mux_v
    port map (
            O => \N__7417\,
            I => \N__7387\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__7408\,
            I => \N__7387\
        );

    \I__1306\ : InMux
    port map (
            O => \N__7407\,
            I => \N__7384\
        );

    \I__1305\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7381\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__7403\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1303\ : Odrv12
    port map (
            O => \N__7400\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__7397\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__7394\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__7387\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__7384\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__7381\,
            I => \U409_AUTOCONFIG.BRIDGE_CONFZ0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__7366\,
            I => \N__7363\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7363\,
            I => \U409_CIA.un1_CIA_CLK_COUNT_3_2\
        );

    \I__1295\ : InMux
    port map (
            O => \N__7360\,
            I => \N__7354\
        );

    \I__1294\ : InMux
    port map (
            O => \N__7359\,
            I => \N__7351\
        );

    \I__1293\ : InMux
    port map (
            O => \N__7358\,
            I => \N__7346\
        );

    \I__1292\ : InMux
    port map (
            O => \N__7357\,
            I => \N__7346\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__7354\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__7351\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7346\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_2\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__7339\,
            I => \N__7333\
        );

    \I__1287\ : InMux
    port map (
            O => \N__7338\,
            I => \N__7330\
        );

    \I__1286\ : InMux
    port map (
            O => \N__7337\,
            I => \N__7327\
        );

    \I__1285\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7324\
        );

    \I__1284\ : InMux
    port map (
            O => \N__7333\,
            I => \N__7321\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__7330\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__7327\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__7324\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__7321\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_5\
        );

    \I__1279\ : CascadeMux
    port map (
            O => \N__7312\,
            I => \N__7308\
        );

    \I__1278\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7303\
        );

    \I__1277\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7300\
        );

    \I__1276\ : InMux
    port map (
            O => \N__7307\,
            I => \N__7297\
        );

    \I__1275\ : InMux
    port map (
            O => \N__7306\,
            I => \N__7294\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__7303\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__7300\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__7297\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__7294\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_3\
        );

    \I__1270\ : InMux
    port map (
            O => \N__7285\,
            I => \N__7279\
        );

    \I__1269\ : InMux
    port map (
            O => \N__7284\,
            I => \N__7276\
        );

    \I__1268\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7271\
        );

    \I__1267\ : InMux
    port map (
            O => \N__7282\,
            I => \N__7271\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__7279\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__7276\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__7271\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_4\
        );

    \I__1263\ : CascadeMux
    port map (
            O => \N__7264\,
            I => \U409_CIA.CIA_CLK_COUNT11_3_cascade_\
        );

    \I__1262\ : InMux
    port map (
            O => \N__7261\,
            I => \N__7255\
        );

    \I__1261\ : InMux
    port map (
            O => \N__7260\,
            I => \N__7255\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__7255\,
            I => \U409_CIA.CIA_CLK_COUNT11\
        );

    \I__1259\ : InMux
    port map (
            O => \N__7252\,
            I => \N__7242\
        );

    \I__1258\ : InMux
    port map (
            O => \N__7251\,
            I => \N__7242\
        );

    \I__1257\ : InMux
    port map (
            O => \N__7250\,
            I => \N__7233\
        );

    \I__1256\ : InMux
    port map (
            O => \N__7249\,
            I => \N__7233\
        );

    \I__1255\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7233\
        );

    \I__1254\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7233\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__7242\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__7233\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_0\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__7228\,
            I => \N__7221\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__7227\,
            I => \N__7218\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__7226\,
            I => \N__7215\
        );

    \I__1248\ : InMux
    port map (
            O => \N__7225\,
            I => \N__7211\
        );

    \I__1247\ : InMux
    port map (
            O => \N__7224\,
            I => \N__7206\
        );

    \I__1246\ : InMux
    port map (
            O => \N__7221\,
            I => \N__7206\
        );

    \I__1245\ : InMux
    port map (
            O => \N__7218\,
            I => \N__7199\
        );

    \I__1244\ : InMux
    port map (
            O => \N__7215\,
            I => \N__7199\
        );

    \I__1243\ : InMux
    port map (
            O => \N__7214\,
            I => \N__7199\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__7211\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__7206\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__7199\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_1\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__7192\,
            I => \N__7188\
        );

    \I__1238\ : InMux
    port map (
            O => \N__7191\,
            I => \N__7182\
        );

    \I__1237\ : InMux
    port map (
            O => \N__7188\,
            I => \N__7182\
        );

    \I__1236\ : InMux
    port map (
            O => \N__7187\,
            I => \N__7179\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__7182\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1234\ : LocalMux
    port map (
            O => \N__7179\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_7\
        );

    \I__1233\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7167\
        );

    \I__1232\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7167\
        );

    \I__1231\ : InMux
    port map (
            O => \N__7172\,
            I => \N__7164\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__7167\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1229\ : LocalMux
    port map (
            O => \N__7164\,
            I => \U409_CIA.CIA_CLK_COUNTZ0Z_6\
        );

    \I__1228\ : InMux
    port map (
            O => \N__7159\,
            I => \N__7155\
        );

    \I__1227\ : InMux
    port map (
            O => \N__7158\,
            I => \N__7152\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__7155\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__7152\,
            I => \U409_CIA.CLK_CIA6_4\
        );

    \I__1224\ : CascadeMux
    port map (
            O => \N__7147\,
            I => \U409_ADDRESS_DECODE.N_77_mux_cascade_\
        );

    \I__1223\ : IoInMux
    port map (
            O => \N__7144\,
            I => \N__7141\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__7141\,
            I => \N__7138\
        );

    \I__1221\ : IoSpan4Mux
    port map (
            O => \N__7138\,
            I => \N__7135\
        );

    \I__1220\ : Span4Mux_s3_h
    port map (
            O => \N__7135\,
            I => \N__7132\
        );

    \I__1219\ : Sp12to4
    port map (
            O => \N__7132\,
            I => \N__7129\
        );

    \I__1218\ : Span12Mux_s8_h
    port map (
            O => \N__7129\,
            I => \N__7126\
        );

    \I__1217\ : Odrv12
    port map (
            O => \N__7126\,
            I => \N_22_0_i\
        );

    \I__1216\ : InMux
    port map (
            O => \N__7123\,
            I => \N__7120\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7117\
        );

    \I__1214\ : Span4Mux_h
    port map (
            O => \N__7117\,
            I => \N__7113\
        );

    \I__1213\ : InMux
    port map (
            O => \N__7116\,
            I => \N__7110\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__7113\,
            I => \N__7107\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__7110\,
            I => \N__7104\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__7107\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1209\ : Odrv4
    port map (
            O => \N__7104\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn\
        );

    \I__1208\ : InMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__7093\,
            I => \N__7090\
        );

    \I__1205\ : Span4Mux_v
    port map (
            O => \N__7090\,
            I => \N__7087\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__7087\,
            I => \U409_ADDRESS_DECODE.PORTSIZE_2\
        );

    \I__1203\ : InMux
    port map (
            O => \N__7084\,
            I => \N__7078\
        );

    \I__1202\ : InMux
    port map (
            O => \N__7083\,
            I => \N__7078\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__7078\,
            I => \BRIDGE_BASE_7\
        );

    \I__1200\ : InMux
    port map (
            O => \N__7075\,
            I => \N__7070\
        );

    \I__1199\ : InMux
    port map (
            O => \N__7074\,
            I => \N__7066\
        );

    \I__1198\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7063\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__7070\,
            I => \N__7060\
        );

    \I__1196\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7057\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__7066\,
            I => \N__7052\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__7063\,
            I => \N__7052\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__7060\,
            I => \N__7049\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7046\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__7052\,
            I => \N__7041\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__7049\,
            I => \N__7036\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__7046\,
            I => \N__7036\
        );

    \I__1188\ : InMux
    port map (
            O => \N__7045\,
            I => \N__7033\
        );

    \I__1187\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7030\
        );

    \I__1186\ : Sp12to4
    port map (
            O => \N__7041\,
            I => \N__7021\
        );

    \I__1185\ : Sp12to4
    port map (
            O => \N__7036\,
            I => \N__7021\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__7033\,
            I => \N__7021\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__7030\,
            I => \N__7021\
        );

    \I__1182\ : Odrv12
    port map (
            O => \N__7021\,
            I => \A_c_7\
        );

    \I__1181\ : InMux
    port map (
            O => \N__7018\,
            I => \N__7013\
        );

    \I__1180\ : InMux
    port map (
            O => \N__7017\,
            I => \N__7010\
        );

    \I__1179\ : InMux
    port map (
            O => \N__7016\,
            I => \N__7007\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__7013\,
            I => \N__7004\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__7010\,
            I => \N__6998\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__6998\
        );

    \I__1175\ : Span4Mux_v
    port map (
            O => \N__7004\,
            I => \N__6994\
        );

    \I__1174\ : InMux
    port map (
            O => \N__7003\,
            I => \N__6991\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__6998\,
            I => \N__6988\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6997\,
            I => \N__6985\
        );

    \I__1171\ : Sp12to4
    port map (
            O => \N__6994\,
            I => \N__6976\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__6991\,
            I => \N__6976\
        );

    \I__1169\ : Sp12to4
    port map (
            O => \N__6988\,
            I => \N__6976\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__6985\,
            I => \N__6976\
        );

    \I__1167\ : Span12Mux_h
    port map (
            O => \N__6976\,
            I => \N__6973\
        );

    \I__1166\ : Odrv12
    port map (
            O => \N__6973\,
            I => \A_c_5\
        );

    \I__1165\ : CascadeMux
    port map (
            O => \N__6970\,
            I => \N__6967\
        );

    \I__1164\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6964\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__6964\,
            I => \N__6961\
        );

    \I__1162\ : Span4Mux_h
    port map (
            O => \N__6961\,
            I => \N__6958\
        );

    \I__1161\ : Odrv4
    port map (
            O => \N__6958\,
            I => \U409_AUTOCONFIG.un1_STATE_6Z0Z_1\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6950\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6954\,
            I => \N__6945\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6953\,
            I => \N__6945\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__6950\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6945\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6940\,
            I => \N__6935\
        );

    \I__1154\ : CascadeMux
    port map (
            O => \N__6939\,
            I => \N__6929\
        );

    \I__1153\ : CascadeMux
    port map (
            O => \N__6938\,
            I => \N__6924\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6916\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6916\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__6933\,
            I => \N__6913\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6904\
        );

    \I__1148\ : InMux
    port map (
            O => \N__6929\,
            I => \N__6904\
        );

    \I__1147\ : InMux
    port map (
            O => \N__6928\,
            I => \N__6904\
        );

    \I__1146\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6901\
        );

    \I__1145\ : InMux
    port map (
            O => \N__6924\,
            I => \N__6895\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6923\,
            I => \N__6895\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__6922\,
            I => \N__6891\
        );

    \I__1142\ : CascadeMux
    port map (
            O => \N__6921\,
            I => \N__6888\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__6916\,
            I => \N__6882\
        );

    \I__1140\ : InMux
    port map (
            O => \N__6913\,
            I => \N__6879\
        );

    \I__1139\ : InMux
    port map (
            O => \N__6912\,
            I => \N__6876\
        );

    \I__1138\ : InMux
    port map (
            O => \N__6911\,
            I => \N__6873\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__6904\,
            I => \N__6868\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6901\,
            I => \N__6868\
        );

    \I__1135\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6865\
        );

    \I__1134\ : LocalMux
    port map (
            O => \N__6895\,
            I => \N__6861\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6894\,
            I => \N__6854\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6891\,
            I => \N__6854\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6888\,
            I => \N__6854\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__6887\,
            I => \N__6851\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__6886\,
            I => \N__6846\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__6885\,
            I => \N__6843\
        );

    \I__1127\ : Span4Mux_v
    port map (
            O => \N__6882\,
            I => \N__6838\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__6879\,
            I => \N__6838\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__6876\,
            I => \N__6835\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__6873\,
            I => \N__6832\
        );

    \I__1123\ : Span4Mux_v
    port map (
            O => \N__6868\,
            I => \N__6829\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6865\,
            I => \N__6826\
        );

    \I__1121\ : InMux
    port map (
            O => \N__6864\,
            I => \N__6823\
        );

    \I__1120\ : Span4Mux_v
    port map (
            O => \N__6861\,
            I => \N__6818\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__6854\,
            I => \N__6818\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6851\,
            I => \N__6813\
        );

    \I__1117\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6813\
        );

    \I__1116\ : InMux
    port map (
            O => \N__6849\,
            I => \N__6806\
        );

    \I__1115\ : InMux
    port map (
            O => \N__6846\,
            I => \N__6806\
        );

    \I__1114\ : InMux
    port map (
            O => \N__6843\,
            I => \N__6806\
        );

    \I__1113\ : Span4Mux_v
    port map (
            O => \N__6838\,
            I => \N__6803\
        );

    \I__1112\ : Span4Mux_v
    port map (
            O => \N__6835\,
            I => \N__6798\
        );

    \I__1111\ : Span4Mux_v
    port map (
            O => \N__6832\,
            I => \N__6798\
        );

    \I__1110\ : Span4Mux_h
    port map (
            O => \N__6829\,
            I => \N__6793\
        );

    \I__1109\ : Span4Mux_v
    port map (
            O => \N__6826\,
            I => \N__6793\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6784\
        );

    \I__1107\ : Sp12to4
    port map (
            O => \N__6818\,
            I => \N__6784\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__6813\,
            I => \N__6784\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__6806\,
            I => \N__6784\
        );

    \I__1104\ : Sp12to4
    port map (
            O => \N__6803\,
            I => \N__6779\
        );

    \I__1103\ : Sp12to4
    port map (
            O => \N__6798\,
            I => \N__6779\
        );

    \I__1102\ : Span4Mux_h
    port map (
            O => \N__6793\,
            I => \N__6776\
        );

    \I__1101\ : Span12Mux_h
    port map (
            O => \N__6784\,
            I => \N__6773\
        );

    \I__1100\ : Span12Mux_h
    port map (
            O => \N__6779\,
            I => \N__6768\
        );

    \I__1099\ : Sp12to4
    port map (
            O => \N__6776\,
            I => \N__6768\
        );

    \I__1098\ : Span12Mux_v
    port map (
            O => \N__6773\,
            I => \N__6765\
        );

    \I__1097\ : Span12Mux_v
    port map (
            O => \N__6768\,
            I => \N__6762\
        );

    \I__1096\ : Odrv12
    port map (
            O => \N__6765\,
            I => \A_c_1\
        );

    \I__1095\ : Odrv12
    port map (
            O => \N__6762\,
            I => \A_c_1\
        );

    \I__1094\ : CascadeMux
    port map (
            O => \N__6757\,
            I => \U409_AUTOCONFIG.un1_STATE_6_0_cascade_\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__6754\,
            I => \N__6749\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6746\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__6752\,
            I => \N__6741\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6749\,
            I => \N__6738\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__6746\,
            I => \N__6735\
        );

    \I__1088\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6728\
        );

    \I__1087\ : InMux
    port map (
            O => \N__6744\,
            I => \N__6728\
        );

    \I__1086\ : InMux
    port map (
            O => \N__6741\,
            I => \N__6728\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6738\,
            I => \N__6725\
        );

    \I__1084\ : Span4Mux_h
    port map (
            O => \N__6735\,
            I => \N__6722\
        );

    \I__1083\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6719\
        );

    \I__1082\ : Span4Mux_v
    port map (
            O => \N__6725\,
            I => \N__6716\
        );

    \I__1081\ : Span4Mux_v
    port map (
            O => \N__6722\,
            I => \N__6713\
        );

    \I__1080\ : Span4Mux_h
    port map (
            O => \N__6719\,
            I => \N__6710\
        );

    \I__1079\ : Sp12to4
    port map (
            O => \N__6716\,
            I => \N__6707\
        );

    \I__1078\ : Sp12to4
    port map (
            O => \N__6713\,
            I => \N__6702\
        );

    \I__1077\ : Sp12to4
    port map (
            O => \N__6710\,
            I => \N__6702\
        );

    \I__1076\ : Span12Mux_h
    port map (
            O => \N__6707\,
            I => \N__6699\
        );

    \I__1075\ : Span12Mux_v
    port map (
            O => \N__6702\,
            I => \N__6696\
        );

    \I__1074\ : Odrv12
    port map (
            O => \N__6699\,
            I => \D_in_6\
        );

    \I__1073\ : Odrv12
    port map (
            O => \N__6696\,
            I => \D_in_6\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6691\,
            I => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_\
        );

    \I__1071\ : CascadeMux
    port map (
            O => \N__6688\,
            I => \N__6685\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6684\,
            I => \N__6679\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6679\,
            I => \BRIDGE_BASE_6\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6676\,
            I => \N__6673\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__6673\,
            I => \N__6669\
        );

    \I__1065\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6666\
        );

    \I__1064\ : Span4Mux_h
    port map (
            O => \N__6669\,
            I => \N__6661\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__6666\,
            I => \N__6661\
        );

    \I__1062\ : Odrv4
    port map (
            O => \N__6661\,
            I => \CIA_SPACE\
        );

    \I__1061\ : CascadeMux
    port map (
            O => \N__6658\,
            I => \U409_CIA.VMA_RNOZ0Z_0_cascade_\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6655\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\
        );

    \I__1059\ : IoInMux
    port map (
            O => \N__6652\,
            I => \N__6649\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6649\,
            I => \N__6646\
        );

    \I__1057\ : IoSpan4Mux
    port map (
            O => \N__6646\,
            I => \N__6643\
        );

    \I__1056\ : Span4Mux_s2_v
    port map (
            O => \N__6643\,
            I => \N__6640\
        );

    \I__1055\ : Span4Mux_h
    port map (
            O => \N__6640\,
            I => \N__6637\
        );

    \I__1054\ : Sp12to4
    port map (
            O => \N__6637\,
            I => \N__6634\
        );

    \I__1053\ : Span12Mux_v
    port map (
            O => \N__6634\,
            I => \N__6631\
        );

    \I__1052\ : Odrv12
    port map (
            O => \N__6631\,
            I => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__6625\,
            I => \N__6621\
        );

    \I__1049\ : InMux
    port map (
            O => \N__6624\,
            I => \N__6618\
        );

    \I__1048\ : Span4Mux_h
    port map (
            O => \N__6621\,
            I => \N__6614\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6618\,
            I => \N__6611\
        );

    \I__1046\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6608\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6614\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__6611\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6608\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\
        );

    \I__1042\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__1041\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6595\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__6595\,
            I => \BRIDGE_BASE_0\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6592\,
            I => \N__6589\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6586\
        );

    \I__1037\ : Odrv4
    port map (
            O => \N__6586\,
            I => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4\
        );

    \I__1036\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6580\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__6580\,
            I => \N__6577\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__6577\,
            I => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3\
        );

    \I__1033\ : CascadeMux
    port map (
            O => \N__6574\,
            I => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_\
        );

    \I__1032\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6568\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__6568\,
            I => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2\
        );

    \I__1030\ : IoInMux
    port map (
            O => \N__6565\,
            I => \N__6562\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__6562\,
            I => \N__6559\
        );

    \I__1028\ : IoSpan4Mux
    port map (
            O => \N__6559\,
            I => \N__6556\
        );

    \I__1027\ : Sp12to4
    port map (
            O => \N__6556\,
            I => \N__6553\
        );

    \I__1026\ : Span12Mux_s7_h
    port map (
            O => \N__6553\,
            I => \N__6550\
        );

    \I__1025\ : Span12Mux_h
    port map (
            O => \N__6550\,
            I => \N__6547\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__6547\,
            I => \U409_ADDRESS_DECODE_un1_BREG_ENn_i\
        );

    \I__1023\ : InMux
    port map (
            O => \N__6544\,
            I => \N__6540\
        );

    \I__1022\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6536\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__6540\,
            I => \N__6530\
        );

    \I__1020\ : InMux
    port map (
            O => \N__6539\,
            I => \N__6527\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__6536\,
            I => \N__6524\
        );

    \I__1018\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6519\
        );

    \I__1017\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6519\
        );

    \I__1016\ : InMux
    port map (
            O => \N__6533\,
            I => \N__6515\
        );

    \I__1015\ : Span4Mux_v
    port map (
            O => \N__6530\,
            I => \N__6506\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__6527\,
            I => \N__6506\
        );

    \I__1013\ : Span4Mux_h
    port map (
            O => \N__6524\,
            I => \N__6506\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__6519\,
            I => \N__6506\
        );

    \I__1011\ : InMux
    port map (
            O => \N__6518\,
            I => \N__6503\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__6515\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__6506\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6503\,
            I => \U409_AUTOCONFIG.LIDE_CONFZ0\
        );

    \I__1007\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6493\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6490\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__6490\,
            I => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0\
        );

    \I__1004\ : InMux
    port map (
            O => \N__6487\,
            I => \N__6484\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6484\,
            I => \N__6480\
        );

    \I__1002\ : InMux
    port map (
            O => \N__6483\,
            I => \N__6477\
        );

    \I__1001\ : Odrv4
    port map (
            O => \N__6480\,
            I => \BRIDGE_BASE_4\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__6477\,
            I => \BRIDGE_BASE_4\
        );

    \I__999\ : InMux
    port map (
            O => \N__6472\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\
        );

    \I__998\ : InMux
    port map (
            O => \N__6469\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\
        );

    \I__997\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6463\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6463\,
            I => \U409_CIA.CLK_CIA6_3\
        );

    \I__995\ : InMux
    port map (
            O => \N__6460\,
            I => \N__6457\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__6457\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\
        );

    \I__993\ : IoInMux
    port map (
            O => \N__6454\,
            I => \N__6451\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__6451\,
            I => \N__6448\
        );

    \I__991\ : IoSpan4Mux
    port map (
            O => \N__6448\,
            I => \N__6445\
        );

    \I__990\ : Sp12to4
    port map (
            O => \N__6445\,
            I => \N__6442\
        );

    \I__989\ : Span12Mux_s7_h
    port map (
            O => \N__6442\,
            I => \N__6439\
        );

    \I__988\ : Span12Mux_h
    port map (
            O => \N__6439\,
            I => \N__6436\
        );

    \I__987\ : Odrv12
    port map (
            O => \N__6436\,
            I => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\
        );

    \I__986\ : CascadeMux
    port map (
            O => \N__6433\,
            I => \N__6430\
        );

    \I__985\ : InMux
    port map (
            O => \N__6430\,
            I => \N__6426\
        );

    \I__984\ : InMux
    port map (
            O => \N__6429\,
            I => \N__6423\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__6426\,
            I => \BRIDGE_BASE_2\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__6423\,
            I => \BRIDGE_BASE_2\
        );

    \I__981\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6415\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__6415\,
            I => \U409_AUTOCONFIG.AC_STARTZ0\
        );

    \I__979\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6409\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__6409\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__6406\,
            I => \U409_CIA.CLK_CIA_r_1_0_cascade_\
        );

    \I__976\ : InMux
    port map (
            O => \N__6403\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\
        );

    \I__975\ : InMux
    port map (
            O => \N__6400\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\
        );

    \I__974\ : InMux
    port map (
            O => \N__6397\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\
        );

    \I__973\ : InMux
    port map (
            O => \N__6394\,
            I => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\
        );

    \I__972\ : InMux
    port map (
            O => \N__6391\,
            I => \N__6388\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__6388\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_0\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__6385\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_\
        );

    \I__969\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6375\
        );

    \I__968\ : InMux
    port map (
            O => \N__6381\,
            I => \N__6375\
        );

    \I__967\ : InMux
    port map (
            O => \N__6380\,
            I => \N__6372\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__6375\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__6372\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0\
        );

    \I__964\ : IoInMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6361\
        );

    \I__962\ : IoSpan4Mux
    port map (
            O => \N__6361\,
            I => \N__6358\
        );

    \I__961\ : Sp12to4
    port map (
            O => \N__6358\,
            I => \N__6355\
        );

    \I__960\ : Span12Mux_s7_v
    port map (
            O => \N__6355\,
            I => \N__6352\
        );

    \I__959\ : Odrv12
    port map (
            O => \N__6352\,
            I => \D_OUT_0\
        );

    \I__958\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6345\
        );

    \I__957\ : InMux
    port map (
            O => \N__6348\,
            I => \N__6342\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__6345\,
            I => \U409_AUTOCONFIG.N_90\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__6342\,
            I => \U409_AUTOCONFIG.N_90\
        );

    \I__954\ : InMux
    port map (
            O => \N__6337\,
            I => \N__6334\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__6334\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\
        );

    \I__952\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6328\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__6328\,
            I => \U409_AUTOCONFIG.N_98\
        );

    \I__950\ : InMux
    port map (
            O => \N__6325\,
            I => \N__6322\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__6322\,
            I => \N__6319\
        );

    \I__948\ : Span12Mux_h
    port map (
            O => \N__6319\,
            I => \N__6316\
        );

    \I__947\ : Span12Mux_v
    port map (
            O => \N__6316\,
            I => \N__6313\
        );

    \I__946\ : Odrv12
    port map (
            O => \N__6313\,
            I => \CPUCONFn_c\
        );

    \I__945\ : CascadeMux
    port map (
            O => \N__6310\,
            I => \U409_AUTOCONFIG.STATE4_cascade_\
        );

    \I__944\ : InMux
    port map (
            O => \N__6307\,
            I => \N__6303\
        );

    \I__943\ : InMux
    port map (
            O => \N__6306\,
            I => \N__6300\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6295\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__6300\,
            I => \N__6295\
        );

    \I__940\ : Span4Mux_v
    port map (
            O => \N__6295\,
            I => \N__6292\
        );

    \I__939\ : Odrv4
    port map (
            O => \N__6292\,
            I => \U409_AUTOCONFIG.N_104\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__6289\,
            I => \U409_AUTOCONFIG.N_103_cascade_\
        );

    \I__937\ : InMux
    port map (
            O => \N__6286\,
            I => \N__6283\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__6283\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\
        );

    \I__935\ : CEMux
    port map (
            O => \N__6280\,
            I => \N__6275\
        );

    \I__934\ : CEMux
    port map (
            O => \N__6279\,
            I => \N__6272\
        );

    \I__933\ : CEMux
    port map (
            O => \N__6278\,
            I => \N__6269\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6264\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6272\,
            I => \N__6261\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__6269\,
            I => \N__6258\
        );

    \I__929\ : CEMux
    port map (
            O => \N__6268\,
            I => \N__6255\
        );

    \I__928\ : CEMux
    port map (
            O => \N__6267\,
            I => \N__6252\
        );

    \I__927\ : Span4Mux_v
    port map (
            O => \N__6264\,
            I => \N__6249\
        );

    \I__926\ : Span4Mux_h
    port map (
            O => \N__6261\,
            I => \N__6246\
        );

    \I__925\ : Span4Mux_h
    port map (
            O => \N__6258\,
            I => \N__6243\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6255\,
            I => \N__6240\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__6252\,
            I => \N__6237\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__6249\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__6246\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__920\ : Odrv4
    port map (
            O => \N__6243\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__919\ : Odrv4
    port map (
            O => \N__6240\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__918\ : Odrv4
    port map (
            O => \N__6237\,
            I => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\
        );

    \I__917\ : InMux
    port map (
            O => \N__6226\,
            I => \N__6205\
        );

    \I__916\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6205\
        );

    \I__915\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6202\
        );

    \I__914\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6199\
        );

    \I__913\ : InMux
    port map (
            O => \N__6222\,
            I => \N__6196\
        );

    \I__912\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6187\
        );

    \I__911\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6187\
        );

    \I__910\ : InMux
    port map (
            O => \N__6219\,
            I => \N__6187\
        );

    \I__909\ : InMux
    port map (
            O => \N__6218\,
            I => \N__6187\
        );

    \I__908\ : InMux
    port map (
            O => \N__6217\,
            I => \N__6182\
        );

    \I__907\ : InMux
    port map (
            O => \N__6216\,
            I => \N__6182\
        );

    \I__906\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6177\
        );

    \I__905\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6177\
        );

    \I__904\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6174\
        );

    \I__903\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6169\
        );

    \I__902\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6169\
        );

    \I__901\ : InMux
    port map (
            O => \N__6210\,
            I => \N__6166\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__6205\,
            I => \N__6161\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__6202\,
            I => \N__6161\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__6199\,
            I => \N__6156\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6156\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6143\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6143\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__6177\,
            I => \N__6143\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6143\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6143\
        );

    \I__891\ : LocalMux
    port map (
            O => \N__6166\,
            I => \N__6143\
        );

    \I__890\ : Span4Mux_v
    port map (
            O => \N__6161\,
            I => \N__6139\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__6156\,
            I => \N__6136\
        );

    \I__888\ : Span4Mux_v
    port map (
            O => \N__6143\,
            I => \N__6133\
        );

    \I__887\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6130\
        );

    \I__886\ : Sp12to4
    port map (
            O => \N__6139\,
            I => \N__6121\
        );

    \I__885\ : Sp12to4
    port map (
            O => \N__6136\,
            I => \N__6121\
        );

    \I__884\ : Sp12to4
    port map (
            O => \N__6133\,
            I => \N__6121\
        );

    \I__883\ : LocalMux
    port map (
            O => \N__6130\,
            I => \N__6121\
        );

    \I__882\ : Odrv12
    port map (
            O => \N__6121\,
            I => \A_c_4\
        );

    \I__881\ : CascadeMux
    port map (
            O => \N__6118\,
            I => \N__6113\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__6117\,
            I => \N__6107\
        );

    \I__879\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6100\
        );

    \I__878\ : InMux
    port map (
            O => \N__6113\,
            I => \N__6100\
        );

    \I__877\ : InMux
    port map (
            O => \N__6112\,
            I => \N__6095\
        );

    \I__876\ : InMux
    port map (
            O => \N__6111\,
            I => \N__6095\
        );

    \I__875\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6092\
        );

    \I__874\ : InMux
    port map (
            O => \N__6107\,
            I => \N__6088\
        );

    \I__873\ : InMux
    port map (
            O => \N__6106\,
            I => \N__6085\
        );

    \I__872\ : CascadeMux
    port map (
            O => \N__6105\,
            I => \N__6081\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__6100\,
            I => \N__6073\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__6095\,
            I => \N__6073\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__6092\,
            I => \N__6073\
        );

    \I__868\ : InMux
    port map (
            O => \N__6091\,
            I => \N__6070\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__6088\,
            I => \N__6067\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__6085\,
            I => \N__6064\
        );

    \I__865\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6061\
        );

    \I__864\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6058\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__6080\,
            I => \N__6055\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__6073\,
            I => \N__6052\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__6070\,
            I => \N__6046\
        );

    \I__860\ : Span4Mux_h
    port map (
            O => \N__6067\,
            I => \N__6036\
        );

    \I__859\ : Span4Mux_v
    port map (
            O => \N__6064\,
            I => \N__6036\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6036\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__6058\,
            I => \N__6036\
        );

    \I__856\ : InMux
    port map (
            O => \N__6055\,
            I => \N__6033\
        );

    \I__855\ : Span4Mux_h
    port map (
            O => \N__6052\,
            I => \N__6030\
        );

    \I__854\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6023\
        );

    \I__853\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6023\
        );

    \I__852\ : InMux
    port map (
            O => \N__6049\,
            I => \N__6023\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__6046\,
            I => \N__6020\
        );

    \I__850\ : InMux
    port map (
            O => \N__6045\,
            I => \N__6017\
        );

    \I__849\ : Span4Mux_v
    port map (
            O => \N__6036\,
            I => \N__6014\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__6033\,
            I => \N__6011\
        );

    \I__847\ : Sp12to4
    port map (
            O => \N__6030\,
            I => \N__6002\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__6023\,
            I => \N__6002\
        );

    \I__845\ : Sp12to4
    port map (
            O => \N__6020\,
            I => \N__6002\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__6002\
        );

    \I__843\ : Span4Mux_h
    port map (
            O => \N__6014\,
            I => \N__5997\
        );

    \I__842\ : Span4Mux_v
    port map (
            O => \N__6011\,
            I => \N__5997\
        );

    \I__841\ : Span12Mux_h
    port map (
            O => \N__6002\,
            I => \N__5994\
        );

    \I__840\ : Span4Mux_h
    port map (
            O => \N__5997\,
            I => \N__5991\
        );

    \I__839\ : Span12Mux_v
    port map (
            O => \N__5994\,
            I => \N__5988\
        );

    \I__838\ : Sp12to4
    port map (
            O => \N__5991\,
            I => \N__5985\
        );

    \I__837\ : Odrv12
    port map (
            O => \N__5988\,
            I => \A_c_2\
        );

    \I__836\ : Odrv12
    port map (
            O => \N__5985\,
            I => \A_c_2\
        );

    \I__835\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5972\
        );

    \I__834\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5972\
        );

    \I__833\ : InMux
    port map (
            O => \N__5978\,
            I => \N__5969\
        );

    \I__832\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5965\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5957\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5969\,
            I => \N__5954\
        );

    \I__829\ : InMux
    port map (
            O => \N__5968\,
            I => \N__5951\
        );

    \I__828\ : InMux
    port map (
            O => \N__5965\,
            I => \N__5947\
        );

    \I__827\ : InMux
    port map (
            O => \N__5964\,
            I => \N__5940\
        );

    \I__826\ : InMux
    port map (
            O => \N__5963\,
            I => \N__5940\
        );

    \I__825\ : InMux
    port map (
            O => \N__5962\,
            I => \N__5940\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__5961\,
            I => \N__5936\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__5960\,
            I => \N__5932\
        );

    \I__822\ : Span4Mux_v
    port map (
            O => \N__5957\,
            I => \N__5928\
        );

    \I__821\ : Span4Mux_v
    port map (
            O => \N__5954\,
            I => \N__5925\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__5951\,
            I => \N__5922\
        );

    \I__819\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5919\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__5947\,
            I => \N__5914\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5914\
        );

    \I__816\ : InMux
    port map (
            O => \N__5939\,
            I => \N__5911\
        );

    \I__815\ : InMux
    port map (
            O => \N__5936\,
            I => \N__5902\
        );

    \I__814\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5902\
        );

    \I__813\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5902\
        );

    \I__812\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5902\
        );

    \I__811\ : Odrv4
    port map (
            O => \N__5928\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__810\ : Odrv4
    port map (
            O => \N__5925\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__809\ : Odrv4
    port map (
            O => \N__5922\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5919\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__807\ : Odrv4
    port map (
            O => \N__5914\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__5911\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__5902\,
            I => \U409_AUTOCONFIG.N_109\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__5887\,
            I => \N__5883\
        );

    \I__803\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5878\
        );

    \I__802\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5878\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__5878\,
            I => \N__5875\
        );

    \I__800\ : Odrv4
    port map (
            O => \N__5875\,
            I => \U409_AUTOCONFIG.N_115\
        );

    \I__799\ : CascadeMux
    port map (
            O => \N__5872\,
            I => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\
        );

    \I__798\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5866\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__5866\,
            I => \N__5862\
        );

    \I__796\ : InMux
    port map (
            O => \N__5865\,
            I => \N__5859\
        );

    \I__795\ : Span4Mux_v
    port map (
            O => \N__5862\,
            I => \N__5856\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__5859\,
            I => \N__5853\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__5856\,
            I => \U409_AUTOCONFIG.N_119\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__5853\,
            I => \U409_AUTOCONFIG.N_119\
        );

    \I__791\ : InMux
    port map (
            O => \N__5848\,
            I => \N__5845\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__5842\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_3\
        );

    \I__788\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \U409_AUTOCONFIG.D_OUT_sm0_0_cascade_\
        );

    \I__787\ : IoInMux
    port map (
            O => \N__5836\,
            I => \N__5833\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__5833\,
            I => \N__5830\
        );

    \I__785\ : Span4Mux_s1_v
    port map (
            O => \N__5830\,
            I => \N__5827\
        );

    \I__784\ : Span4Mux_v
    port map (
            O => \N__5827\,
            I => \N__5824\
        );

    \I__783\ : Span4Mux_v
    port map (
            O => \N__5824\,
            I => \N__5821\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__5821\,
            I => \N__5818\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__5818\,
            I => \D_OUT_3\
        );

    \I__780\ : InMux
    port map (
            O => \N__5815\,
            I => \N__5812\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5812\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\
        );

    \I__778\ : InMux
    port map (
            O => \N__5809\,
            I => \N__5806\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__5806\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\
        );

    \I__776\ : InMux
    port map (
            O => \N__5803\,
            I => \N__5800\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__5800\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\
        );

    \I__774\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__5791\,
            I => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_\
        );

    \I__771\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5785\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__5785\,
            I => \N__5782\
        );

    \I__769\ : Span4Mux_v
    port map (
            O => \N__5782\,
            I => \N__5779\
        );

    \I__768\ : Odrv4
    port map (
            O => \N__5779\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_2\
        );

    \I__767\ : IoInMux
    port map (
            O => \N__5776\,
            I => \N__5773\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5773\,
            I => \N__5770\
        );

    \I__765\ : Span4Mux_s3_v
    port map (
            O => \N__5770\,
            I => \N__5767\
        );

    \I__764\ : Sp12to4
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__763\ : Span12Mux_h
    port map (
            O => \N__5764\,
            I => \N__5761\
        );

    \I__762\ : Span12Mux_v
    port map (
            O => \N__5761\,
            I => \N__5758\
        );

    \I__761\ : Odrv12
    port map (
            O => \N__5758\,
            I => \PORTSIZE_0_i\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5755\,
            I => \N__5751\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__5754\,
            I => \N__5748\
        );

    \I__758\ : InMux
    port map (
            O => \N__5751\,
            I => \N__5744\
        );

    \I__757\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5741\
        );

    \I__756\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5738\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__5744\,
            I => \N__5731\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5731\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5727\
        );

    \I__752\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5724\
        );

    \I__751\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5721\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__5731\,
            I => \N__5718\
        );

    \I__749\ : InMux
    port map (
            O => \N__5730\,
            I => \N__5715\
        );

    \I__748\ : Span4Mux_h
    port map (
            O => \N__5727\,
            I => \N__5708\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__5724\,
            I => \N__5708\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__5721\,
            I => \N__5708\
        );

    \I__745\ : Sp12to4
    port map (
            O => \N__5718\,
            I => \N__5705\
        );

    \I__744\ : LocalMux
    port map (
            O => \N__5715\,
            I => \N__5702\
        );

    \I__743\ : Sp12to4
    port map (
            O => \N__5708\,
            I => \N__5699\
        );

    \I__742\ : Span12Mux_h
    port map (
            O => \N__5705\,
            I => \N__5694\
        );

    \I__741\ : Span12Mux_v
    port map (
            O => \N__5702\,
            I => \N__5694\
        );

    \I__740\ : Span12Mux_v
    port map (
            O => \N__5699\,
            I => \N__5691\
        );

    \I__739\ : Span12Mux_v
    port map (
            O => \N__5694\,
            I => \N__5688\
        );

    \I__738\ : Odrv12
    port map (
            O => \N__5691\,
            I => \A_c_3\
        );

    \I__737\ : Odrv12
    port map (
            O => \N__5688\,
            I => \A_c_3\
        );

    \I__736\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5679\
        );

    \I__735\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5676\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__5679\,
            I => \N__5671\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5676\,
            I => \N__5666\
        );

    \I__732\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5661\
        );

    \I__731\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5661\
        );

    \I__730\ : Span4Mux_v
    port map (
            O => \N__5671\,
            I => \N__5658\
        );

    \I__729\ : InMux
    port map (
            O => \N__5670\,
            I => \N__5655\
        );

    \I__728\ : InMux
    port map (
            O => \N__5669\,
            I => \N__5652\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__5666\,
            I => \N__5649\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__5661\,
            I => \N__5640\
        );

    \I__725\ : Sp12to4
    port map (
            O => \N__5658\,
            I => \N__5640\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5655\,
            I => \N__5640\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5652\,
            I => \N__5640\
        );

    \I__722\ : Span4Mux_h
    port map (
            O => \N__5649\,
            I => \N__5637\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__5640\,
            I => \A_c_6\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__5637\,
            I => \A_c_6\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \U409_AUTOCONFIG.N_109_cascade_\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__5629\,
            I => \N__5625\
        );

    \I__717\ : InMux
    port map (
            O => \N__5628\,
            I => \N__5620\
        );

    \I__716\ : InMux
    port map (
            O => \N__5625\,
            I => \N__5620\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5620\,
            I => \U409_AUTOCONFIG.N_117\
        );

    \I__714\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5614\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__5614\,
            I => \N__5610\
        );

    \I__712\ : InMux
    port map (
            O => \N__5613\,
            I => \N__5607\
        );

    \I__711\ : Odrv12
    port map (
            O => \N__5610\,
            I => \U409_AUTOCONFIG.N_113\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__5607\,
            I => \U409_AUTOCONFIG.N_113\
        );

    \I__709\ : InMux
    port map (
            O => \N__5602\,
            I => \N__5599\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5599\,
            I => \N__5596\
        );

    \I__707\ : Span4Mux_v
    port map (
            O => \N__5596\,
            I => \N__5593\
        );

    \I__706\ : Sp12to4
    port map (
            O => \N__5593\,
            I => \N__5590\
        );

    \I__705\ : Span12Mux_h
    port map (
            O => \N__5590\,
            I => \N__5587\
        );

    \I__704\ : Span12Mux_h
    port map (
            O => \N__5587\,
            I => \N__5584\
        );

    \I__703\ : Span12Mux_v
    port map (
            O => \N__5584\,
            I => \N__5581\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__5581\,
            I => \AUTOBOOT_c\
        );

    \I__701\ : InMux
    port map (
            O => \N__5578\,
            I => \N__5575\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5575\,
            I => \N__5572\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5572\,
            I => \U409_AUTOCONFIG.N_101\
        );

    \I__698\ : InMux
    port map (
            O => \N__5569\,
            I => \N__5566\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5566\,
            I => \U409_AUTOCONFIG.PR_OUTZ0Z_1\
        );

    \I__696\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5560\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__5560\,
            I => \U409_AUTOCONFIG.N_91\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__5557\,
            I => \U409_AUTOCONFIG.N_91_cascade_\
        );

    \I__693\ : InMux
    port map (
            O => \N__5554\,
            I => \N__5551\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__5551\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\
        );

    \I__691\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__690\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5542\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5542\,
            I => \U409_AUTOCONFIG.N_216_3\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5539\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_\
        );

    \I__687\ : InMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__5533\,
            I => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\
        );

    \I__685\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__684\ : LocalMux
    port map (
            O => \N__5527\,
            I => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\
        );

    \I__683\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5521\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5518\
        );

    \I__681\ : Odrv4
    port map (
            O => \N__5518\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\
        );

    \I__680\ : InMux
    port map (
            O => \N__5515\,
            I => \N__5511\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__5514\,
            I => \N__5508\
        );

    \I__678\ : LocalMux
    port map (
            O => \N__5511\,
            I => \N__5505\
        );

    \I__677\ : InMux
    port map (
            O => \N__5508\,
            I => \N__5502\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__5505\,
            I => \U409_AUTOCONFIG.N_116\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5502\,
            I => \U409_AUTOCONFIG.N_116\
        );

    \I__674\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5494\
        );

    \I__673\ : LocalMux
    port map (
            O => \N__5494\,
            I => \N__5489\
        );

    \I__672\ : InMux
    port map (
            O => \N__5493\,
            I => \N__5486\
        );

    \I__671\ : InMux
    port map (
            O => \N__5492\,
            I => \N__5483\
        );

    \I__670\ : Odrv4
    port map (
            O => \N__5489\,
            I => \U409_AUTOCONFIG.N_89\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__5486\,
            I => \U409_AUTOCONFIG.N_89\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__5483\,
            I => \U409_AUTOCONFIG.N_89\
        );

    \I__667\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5473\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__5473\,
            I => \N__5470\
        );

    \I__665\ : Odrv4
    port map (
            O => \N__5470\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_8\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \N__5464\
        );

    \I__663\ : InMux
    port map (
            O => \N__5464\,
            I => \N__5461\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__661\ : Span4Mux_h
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__660\ : Span4Mux_v
    port map (
            O => \N__5455\,
            I => \N__5452\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__5452\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_9\
        );

    \I__658\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5446\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__5446\,
            I => \U409_ADDRESS_DECODE_AUTOVECTOR_10\
        );

    \I__656\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5440\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__5440\,
            I => \U409_AUTOCONFIG.N_99\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__5437\,
            I => \N__5434\
        );

    \I__653\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5431\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__5431\,
            I => \N__5428\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__5428\,
            I => \U409_AUTOCONFIG.N_100\
        );

    \I__650\ : CascadeMux
    port map (
            O => \N__5425\,
            I => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\
        );

    \I__649\ : IoInMux
    port map (
            O => \N__5422\,
            I => \N__5419\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__5419\,
            I => \N__5416\
        );

    \I__647\ : Span4Mux_s2_v
    port map (
            O => \N__5416\,
            I => \N__5413\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__5413\,
            I => \N__5410\
        );

    \I__645\ : Span4Mux_v
    port map (
            O => \N__5410\,
            I => \N__5407\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__5407\,
            I => \D_OUT_2\
        );

    \I__643\ : IoInMux
    port map (
            O => \N__5404\,
            I => \N__5401\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__5401\,
            I => \N__5398\
        );

    \I__641\ : Span4Mux_s1_v
    port map (
            O => \N__5398\,
            I => \N__5395\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__5395\,
            I => \N__5392\
        );

    \I__639\ : Span4Mux_v
    port map (
            O => \N__5392\,
            I => \N__5389\
        );

    \I__638\ : Odrv4
    port map (
            O => \N__5389\,
            I => \D_OUT_1\
        );

    \I__637\ : InMux
    port map (
            O => \N__5386\,
            I => \N__5383\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__5383\,
            I => \U409_AUTOCONFIG.N_111\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__5380\,
            I => \U409_AUTOCONFIG.N_105_cascade_\
        );

    \I__634\ : InMux
    port map (
            O => \N__5377\,
            I => \N__5374\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__5374\,
            I => \N__5370\
        );

    \I__632\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5367\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__5370\,
            I => \PRO_BASE_1\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__5367\,
            I => \PRO_BASE_1\
        );

    \I__629\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_\
        );

    \I__628\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5350\
        );

    \I__627\ : InMux
    port map (
            O => \N__5358\,
            I => \N__5350\
        );

    \I__626\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5350\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__5350\,
            I => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\
        );

    \I__624\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5344\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5341\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__5341\,
            I => \U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__5338\,
            I => \U409_AUTOCONFIG.N_216_3_cascade_\
        );

    \I__620\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5332\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__5332\,
            I => \U409_AUTOCONFIG.N_108\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__5329\,
            I => \U409_AUTOCONFIG.N_108_cascade_\
        );

    \I__617\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5323\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__5323\,
            I => \U409_ADDRESS_DECODE.N_59\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__5320\,
            I => \U409_ADDRESS_DECODE.N_59_cascade_\
        );

    \I__614\ : InMux
    port map (
            O => \N__5317\,
            I => \N__5314\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__5314\,
            I => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\
        );

    \I__612\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5308\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__5308\,
            I => \N__5305\
        );

    \I__610\ : Span4Mux_v
    port map (
            O => \N__5305\,
            I => \N__5301\
        );

    \I__609\ : InMux
    port map (
            O => \N__5304\,
            I => \N__5298\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__5301\,
            I => \N__5293\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__5298\,
            I => \N__5293\
        );

    \I__606\ : Span4Mux_h
    port map (
            O => \N__5293\,
            I => \N__5290\
        );

    \I__605\ : Sp12to4
    port map (
            O => \N__5290\,
            I => \N__5287\
        );

    \I__604\ : Odrv12
    port map (
            O => \N__5287\,
            I => \TT_c_1\
        );

    \I__603\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5281\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__5281\,
            I => \N__5278\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__5278\,
            I => \N__5274\
        );

    \I__600\ : InMux
    port map (
            O => \N__5277\,
            I => \N__5271\
        );

    \I__599\ : Span4Mux_h
    port map (
            O => \N__5274\,
            I => \N__5268\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__5271\,
            I => \N__5265\
        );

    \I__597\ : Sp12to4
    port map (
            O => \N__5268\,
            I => \N__5260\
        );

    \I__596\ : Span12Mux_h
    port map (
            O => \N__5265\,
            I => \N__5260\
        );

    \I__595\ : Odrv12
    port map (
            O => \N__5260\,
            I => \TT_c_0\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \N__5254\
        );

    \I__593\ : InMux
    port map (
            O => \N__5254\,
            I => \N__5251\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__5251\,
            I => \N__5248\
        );

    \I__591\ : Span4Mux_v
    port map (
            O => \N__5248\,
            I => \N__5245\
        );

    \I__590\ : Span4Mux_v
    port map (
            O => \N__5245\,
            I => \N__5242\
        );

    \I__589\ : IoSpan4Mux
    port map (
            O => \N__5242\,
            I => \N__5239\
        );

    \I__588\ : Odrv4
    port map (
            O => \N__5239\,
            I => \TM_c_2\
        );

    \I__587\ : IoInMux
    port map (
            O => \N__5236\,
            I => \N__5233\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__5233\,
            I => \N__5228\
        );

    \I__585\ : IoInMux
    port map (
            O => \N__5232\,
            I => \N__5225\
        );

    \I__584\ : IoInMux
    port map (
            O => \N__5231\,
            I => \N__5222\
        );

    \I__583\ : IoSpan4Mux
    port map (
            O => \N__5228\,
            I => \N__5214\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__5225\,
            I => \N__5214\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__5222\,
            I => \N__5214\
        );

    \I__580\ : IoInMux
    port map (
            O => \N__5221\,
            I => \N__5211\
        );

    \I__579\ : IoSpan4Mux
    port map (
            O => \N__5214\,
            I => \N__5208\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5205\
        );

    \I__577\ : Span4Mux_s3_v
    port map (
            O => \N__5208\,
            I => \N__5200\
        );

    \I__576\ : Span4Mux_s3_v
    port map (
            O => \N__5205\,
            I => \N__5200\
        );

    \I__575\ : Span4Mux_v
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__574\ : Odrv4
    port map (
            O => \N__5197\,
            I => \D_1_i\
        );

    \I__573\ : IoInMux
    port map (
            O => \N__5194\,
            I => \N__5191\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__5191\,
            I => \N__5188\
        );

    \I__571\ : Span4Mux_s1_v
    port map (
            O => \N__5188\,
            I => \N__5185\
        );

    \I__570\ : Sp12to4
    port map (
            O => \N__5185\,
            I => \N__5181\
        );

    \I__569\ : CascadeMux
    port map (
            O => \N__5184\,
            I => \N__5178\
        );

    \I__568\ : Span12Mux_h
    port map (
            O => \N__5181\,
            I => \N__5175\
        );

    \I__567\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5172\
        );

    \I__566\ : Odrv12
    port map (
            O => \N__5175\,
            I => \CONFIGENn_c\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__5172\,
            I => \CONFIGENn_c\
        );

    \I__564\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5163\
        );

    \I__563\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5160\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__5163\,
            I => \PRO_BASE_2\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__5160\,
            I => \PRO_BASE_2\
        );

    \I__560\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5151\
        );

    \I__559\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5148\
        );

    \I__558\ : LocalMux
    port map (
            O => \N__5151\,
            I => \PRO_BASE_0\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__5148\,
            I => \PRO_BASE_0\
        );

    \I__556\ : IoInMux
    port map (
            O => \N__5143\,
            I => \N__5140\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__5140\,
            I => \N__5137\
        );

    \I__554\ : Span4Mux_s0_v
    port map (
            O => \N__5137\,
            I => \N__5134\
        );

    \I__553\ : Sp12to4
    port map (
            O => \N__5134\,
            I => \N__5131\
        );

    \I__552\ : Span12Mux_h
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__551\ : Span12Mux_v
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__550\ : Odrv12
    port map (
            O => \N__5125\,
            I => \U409_ADDRESS_DECODE_un1_BPRO_ENn_i\
        );

    \I__549\ : InMux
    port map (
            O => \N__5122\,
            I => \N__5117\
        );

    \I__548\ : InMux
    port map (
            O => \N__5121\,
            I => \N__5114\
        );

    \I__547\ : InMux
    port map (
            O => \N__5120\,
            I => \N__5111\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__5117\,
            I => \N__5108\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5103\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__5111\,
            I => \N__5103\
        );

    \I__543\ : Sp12to4
    port map (
            O => \N__5108\,
            I => \N__5100\
        );

    \I__542\ : Sp12to4
    port map (
            O => \N__5103\,
            I => \N__5097\
        );

    \I__541\ : Span12Mux_v
    port map (
            O => \N__5100\,
            I => \N__5094\
        );

    \I__540\ : Span12Mux_v
    port map (
            O => \N__5097\,
            I => \N__5091\
        );

    \I__539\ : Odrv12
    port map (
            O => \N__5094\,
            I => \A_c_29\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__5091\,
            I => \A_c_29\
        );

    \I__537\ : CascadeMux
    port map (
            O => \N__5086\,
            I => \U409_ADDRESS_DECODE.N_26_cascade_\
        );

    \I__536\ : InMux
    port map (
            O => \N__5083\,
            I => \N__5080\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__5080\,
            I => \U409_ADDRESS_DECODE.m54Z0Z_1\
        );

    \I__534\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5074\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__5074\,
            I => \N__5071\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__5071\,
            I => \N__5068\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__5068\,
            I => \U409_AUTOCONFIG.un1_A_13Z0Z_3\
        );

    \I__530\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5062\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__5062\,
            I => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0\
        );

    \I__528\ : InMux
    port map (
            O => \N__5059\,
            I => \N__5056\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__5056\,
            I => \N__5052\
        );

    \I__526\ : InMux
    port map (
            O => \N__5055\,
            I => \N__5049\
        );

    \I__525\ : Span4Mux_v
    port map (
            O => \N__5052\,
            I => \N__5044\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__5049\,
            I => \N__5044\
        );

    \I__523\ : Span4Mux_h
    port map (
            O => \N__5044\,
            I => \N__5040\
        );

    \I__522\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5037\
        );

    \I__521\ : Span4Mux_v
    port map (
            O => \N__5040\,
            I => \N__5032\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__5037\,
            I => \N__5032\
        );

    \I__519\ : Span4Mux_h
    port map (
            O => \N__5032\,
            I => \N__5029\
        );

    \I__518\ : Span4Mux_v
    port map (
            O => \N__5029\,
            I => \N__5026\
        );

    \I__517\ : Odrv4
    port map (
            O => \N__5026\,
            I => \A_c_30\
        );

    \I__516\ : InMux
    port map (
            O => \N__5023\,
            I => \N__5019\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__5019\,
            I => \N__5013\
        );

    \I__513\ : InMux
    port map (
            O => \N__5016\,
            I => \N__5009\
        );

    \I__512\ : Span4Mux_h
    port map (
            O => \N__5013\,
            I => \N__5006\
        );

    \I__511\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5003\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__5000\
        );

    \I__509\ : Span4Mux_v
    port map (
            O => \N__5006\,
            I => \N__4995\
        );

    \I__508\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__4995\
        );

    \I__507\ : Span12Mux_h
    port map (
            O => \N__5000\,
            I => \N__4992\
        );

    \I__506\ : Span4Mux_h
    port map (
            O => \N__4995\,
            I => \N__4989\
        );

    \I__505\ : Span12Mux_v
    port map (
            O => \N__4992\,
            I => \N__4986\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__4989\,
            I => \N__4983\
        );

    \I__503\ : Odrv12
    port map (
            O => \N__4986\,
            I => \A_c_31\
        );

    \I__502\ : Odrv4
    port map (
            O => \N__4983\,
            I => \A_c_31\
        );

    \I__501\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4975\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4975\,
            I => \U409_ADDRESS_DECODE.m12Z0Z_5\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__4972\,
            I => \U409_ADDRESS_DECODE.m12Z0Z_0_cascade_\
        );

    \I__498\ : InMux
    port map (
            O => \N__4969\,
            I => \N__4966\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__4966\,
            I => \U409_AUTOCONFIG.un1_A_13Z0Z_1\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__4963\,
            I => \N__4960\
        );

    \I__495\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4956\
        );

    \I__494\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4953\
        );

    \I__493\ : LocalMux
    port map (
            O => \N__4956\,
            I => \N__4950\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__4953\,
            I => \N__4947\
        );

    \I__491\ : Sp12to4
    port map (
            O => \N__4950\,
            I => \N__4944\
        );

    \I__490\ : Span4Mux_v
    port map (
            O => \N__4947\,
            I => \N__4941\
        );

    \I__489\ : Span12Mux_v
    port map (
            O => \N__4944\,
            I => \N__4938\
        );

    \I__488\ : Span4Mux_h
    port map (
            O => \N__4941\,
            I => \N__4935\
        );

    \I__487\ : Odrv12
    port map (
            O => \N__4938\,
            I => \A_c_25\
        );

    \I__486\ : Odrv4
    port map (
            O => \N__4935\,
            I => \A_c_25\
        );

    \I__485\ : CascadeMux
    port map (
            O => \N__4930\,
            I => \N__4927\
        );

    \I__484\ : InMux
    port map (
            O => \N__4927\,
            I => \N__4923\
        );

    \I__483\ : InMux
    port map (
            O => \N__4926\,
            I => \N__4920\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__4923\,
            I => \N__4917\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4920\,
            I => \N__4914\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__4917\,
            I => \N__4911\
        );

    \I__479\ : Sp12to4
    port map (
            O => \N__4914\,
            I => \N__4908\
        );

    \I__478\ : Span4Mux_v
    port map (
            O => \N__4911\,
            I => \N__4905\
        );

    \I__477\ : Span12Mux_v
    port map (
            O => \N__4908\,
            I => \N__4902\
        );

    \I__476\ : Span4Mux_h
    port map (
            O => \N__4905\,
            I => \N__4899\
        );

    \I__475\ : Odrv12
    port map (
            O => \N__4902\,
            I => \A_c_24\
        );

    \I__474\ : Odrv4
    port map (
            O => \N__4899\,
            I => \A_c_24\
        );

    \I__473\ : InMux
    port map (
            O => \N__4894\,
            I => \N__4891\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__4891\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__4888\,
            I => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\
        );

    \I__470\ : InMux
    port map (
            O => \N__4885\,
            I => \N__4879\
        );

    \I__469\ : InMux
    port map (
            O => \N__4884\,
            I => \N__4879\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__4879\,
            I => \N__4876\
        );

    \I__467\ : Span4Mux_v
    port map (
            O => \N__4876\,
            I => \N__4873\
        );

    \I__466\ : Sp12to4
    port map (
            O => \N__4873\,
            I => \N__4870\
        );

    \I__465\ : Odrv12
    port map (
            O => \N__4870\,
            I => \A_c_27\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__4867\,
            I => \N__4863\
        );

    \I__463\ : InMux
    port map (
            O => \N__4866\,
            I => \N__4860\
        );

    \I__462\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4857\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4860\,
            I => \N__4854\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__4857\,
            I => \N__4851\
        );

    \I__459\ : Span4Mux_v
    port map (
            O => \N__4854\,
            I => \N__4846\
        );

    \I__458\ : Span4Mux_v
    port map (
            O => \N__4851\,
            I => \N__4846\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__4846\,
            I => \N__4843\
        );

    \I__456\ : Span4Mux_v
    port map (
            O => \N__4843\,
            I => \N__4840\
        );

    \I__455\ : Span4Mux_h
    port map (
            O => \N__4840\,
            I => \N__4837\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__4837\,
            I => \A_c_28\
        );

    \I__453\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4830\
        );

    \I__452\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4827\
        );

    \I__451\ : LocalMux
    port map (
            O => \N__4830\,
            I => \N__4824\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__4827\,
            I => \N__4821\
        );

    \I__449\ : Span4Mux_v
    port map (
            O => \N__4824\,
            I => \N__4818\
        );

    \I__448\ : Span4Mux_v
    port map (
            O => \N__4821\,
            I => \N__4815\
        );

    \I__447\ : Span4Mux_v
    port map (
            O => \N__4818\,
            I => \N__4812\
        );

    \I__446\ : Span4Mux_v
    port map (
            O => \N__4815\,
            I => \N__4809\
        );

    \I__445\ : Span4Mux_h
    port map (
            O => \N__4812\,
            I => \N__4806\
        );

    \I__444\ : Span4Mux_h
    port map (
            O => \N__4809\,
            I => \N__4803\
        );

    \I__443\ : Odrv4
    port map (
            O => \N__4806\,
            I => \A_c_26\
        );

    \I__442\ : Odrv4
    port map (
            O => \N__4803\,
            I => \A_c_26\
        );

    \I__441\ : IoInMux
    port map (
            O => \N__4798\,
            I => \N__4795\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__4795\,
            I => \N__4792\
        );

    \I__439\ : IoSpan4Mux
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__4789\,
            I => \N__4786\
        );

    \I__437\ : Span12Mux_s1_h
    port map (
            O => \N__4786\,
            I => \N__4783\
        );

    \I__436\ : Span12Mux_v
    port map (
            O => \N__4783\,
            I => \N__4780\
        );

    \I__435\ : Odrv12
    port map (
            O => \N__4780\,
            I => \PPIO_c\
        );

    \I__434\ : IoInMux
    port map (
            O => \N__4777\,
            I => \N__4774\
        );

    \I__433\ : LocalMux
    port map (
            O => \N__4774\,
            I => \N__4771\
        );

    \I__432\ : Span12Mux_s2_h
    port map (
            O => \N__4771\,
            I => \N__4768\
        );

    \I__431\ : Span12Mux_v
    port map (
            O => \N__4768\,
            I => \N__4765\
        );

    \I__430\ : Odrv12
    port map (
            O => \N__4765\,
            I => \SPIO_c\
        );

    \I__429\ : ClkMux
    port map (
            O => \N__4762\,
            I => \N__4723\
        );

    \I__428\ : ClkMux
    port map (
            O => \N__4761\,
            I => \N__4723\
        );

    \I__427\ : ClkMux
    port map (
            O => \N__4760\,
            I => \N__4723\
        );

    \I__426\ : ClkMux
    port map (
            O => \N__4759\,
            I => \N__4723\
        );

    \I__425\ : ClkMux
    port map (
            O => \N__4758\,
            I => \N__4723\
        );

    \I__424\ : ClkMux
    port map (
            O => \N__4757\,
            I => \N__4723\
        );

    \I__423\ : ClkMux
    port map (
            O => \N__4756\,
            I => \N__4723\
        );

    \I__422\ : ClkMux
    port map (
            O => \N__4755\,
            I => \N__4723\
        );

    \I__421\ : ClkMux
    port map (
            O => \N__4754\,
            I => \N__4723\
        );

    \I__420\ : ClkMux
    port map (
            O => \N__4753\,
            I => \N__4723\
        );

    \I__419\ : ClkMux
    port map (
            O => \N__4752\,
            I => \N__4723\
        );

    \I__418\ : ClkMux
    port map (
            O => \N__4751\,
            I => \N__4723\
        );

    \I__417\ : ClkMux
    port map (
            O => \N__4750\,
            I => \N__4723\
        );

    \I__416\ : GlobalMux
    port map (
            O => \N__4723\,
            I => \CLK80_OUT\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            I => \N__4762\
        );

    \INVU409_TRANSFER_ACK.LASTCLK_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            I => \N__4760\
        );

    \INVU409_TRANSFER_ACK.CIA_STATE_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            I => \N__4758\
        );

    \INVU409_TRANSFER_ACK.CIA_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            I => \N__4755\
        );

    \INVU409_TRANSFER_ACK.ROMENnC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            I => \N__4757\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_ENC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            I => \N__4754\
        );

    \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            I => \N__4753\
        );

    \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            I => \N__4751\
        );

    \INVU409_TRANSFER_ACK.TACK_COUNTER_0C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            I => \N__4750\
        );

    \INVU409_AUTOCONFIG.AC_TACKC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            I => \N__11161\
        );

    \INVU409_AUTOCONFIG.STATE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.STATE_1C_net\,
            I => \N__11165\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\,
            I => \N__4752\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            I => \N__4759\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            I => \N__4756\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_5C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            I => \N__11171\
        );

    \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C\ : INV
    port map (
            O => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            I => \N__4761\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_4C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net\,
            I => \N__11170\
        );

    \INVU409_AUTOCONFIG.BRIDGE_BASE_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net\,
            I => \N__11174\
        );

    \INVU409_AUTOCONFIG.LIDE_BASE_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            I => \N__11181\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_2C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            I => \N__11173\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_3C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            I => \N__11180\
        );

    \INVU409_AUTOCONFIG.BRIDGE_OUT_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            I => \N__11172\
        );

    \INVU409_AUTOCONFIG.PR_OUT_1C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.PR_OUT_1C_net\,
            I => \N__11179\
        );

    \INVU409_AUTOCONFIG.LIDE_OUT_0C\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            I => \N__11182\
        );

    \INVU409_AUTOCONFIG.LIDE_CONFC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            I => \N__11183\
        );

    \INVU409_AUTOCONFIG.CONFIGENnC\ : INV
    port map (
            O => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            I => \N__11187\
        );

    \IN_MUX_bfv_14_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_6_0_\
        );

    \IN_MUX_bfv_14_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un3_COUNTER60_1_cry_8\,
            carryinitout => \bfn_14_7_0_\
        );

    \IN_MUX_bfv_17_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_5_0_\
        );

    \IN_MUX_bfv_17_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \U409_TICK.un2_COUNTER50_1_cry_8\,
            carryinitout => \bfn_17_6_0_\
        );

    \IN_MUX_bfv_8_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_12_0_\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__9538\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m12_5_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4885\,
            in1 => \N__5043\,
            in2 => \N__4930\,
            in3 => \N__4866\,
            lcout => \U409_ADDRESS_DECODE.m12Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_9_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__4884\,
            in1 => \N__5120\,
            in2 => \N__4867\,
            in3 => \N__4833\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5682\,
            lcout => \U409_AUTOCONFIG.un1_A_13Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m12_0_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__4834\,
            in1 => \N__11809\,
            in2 => \_gnd_net_\,
            in3 => \N__5121\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.m12Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m12_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5012\,
            in1 => \N__4978\,
            in2 => \N__4972\,
            in3 => \N__4959\,
            lcout => \U409_ADDRESS_DECODE.Z2_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_LC_3_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7735\,
            in1 => \N__9974\,
            in2 => \N__9283\,
            in3 => \N__7805\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m1_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__10174\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9915\,
            lcout => \U409_ADDRESS_DECODE.N_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_3_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__6900\,
            in1 => \N__7044\,
            in2 => \N__6080\,
            in3 => \N__4969\,
            lcout => \U409_AUTOCONFIG.un1_A_13Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_8_LC_3_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9082\,
            in1 => \N__8477\,
            in2 => \N__4963\,
            in3 => \N__4926\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_3_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__7710\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7809\,
            lcout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_4_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9092\,
            in1 => \N__9698\,
            in2 => \N__10018\,
            in3 => \N__10100\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.AUTOCONFIG_SPACEZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOCONFIG_SPACE_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4894\,
            in1 => \N__9375\,
            in2 => \N__4888\,
            in3 => \N__9284\,
            lcout => \AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m13_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9352\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10194\,
            lcout => \U409_ADDRESS_DECODE.CIA_SPACE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BPRO_ENn_i_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110111111111"
        )
    port map (
            in0 => \N__5083\,
            in1 => \N__5167\,
            in2 => \N__5022\,
            in3 => \N__7631\,
            lcout => \U409_ADDRESS_DECODE_un1_BPRO_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m47_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110111011"
        )
    port map (
            in0 => \N__5122\,
            in1 => \N__11876\,
            in2 => \_gnd_net_\,
            in3 => \N__5155\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.N_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m54_1_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000101"
        )
    port map (
            in0 => \N__5059\,
            in1 => \_gnd_net_\,
            in2 => \N__5086\,
            in3 => \N__5377\,
            lcout => \U409_ADDRESS_DECODE.m54Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_13_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__6223\,
            in1 => \N__7017\,
            in2 => \_gnd_net_\,
            in3 => \N__5077\,
            lcout => \U409_AUTOCONFIG.un1_AZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5065\,
            in1 => \N__5747\,
            in2 => \N__5514\,
            in3 => \N__6911\,
            lcout => \U409_AUTOCONFIG.N_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7016\,
            in1 => \N__7045\,
            in2 => \_gnd_net_\,
            in3 => \N__5683\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a4_0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_1_3_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6222\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6091\,
            lcout => \U409_AUTOCONFIG.N_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_10_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5055\,
            in1 => \N__5317\,
            in2 => \_gnd_net_\,
            in3 => \N__5023\,
            lcout => \U409_ADDRESS_DECODE_AUTOVECTOR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_3_0_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__7069\,
            in1 => \N__5669\,
            in2 => \_gnd_net_\,
            in3 => \N__5736\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_7_i_a4_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CIA_SPACE_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__9867\,
            in1 => \N__5326\,
            in2 => \N__8495\,
            in3 => \N__8542\,
            lcout => \CIA_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m3_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9683\,
            in2 => \_gnd_net_\,
            in3 => \N__10045\,
            lcout => \U409_ADDRESS_DECODE.N_59\,
            ltout => \U409_ADDRESS_DECODE.N_59_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.AUTOVECTOR_7_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5311\,
            in1 => \N__5284\,
            in2 => \N__5320\,
            in3 => \N__11883\,
            lcout => \U409_ADDRESS_DECODE.AUTOVECTORZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m41_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__5304\,
            in1 => \N__5277\,
            in2 => \N__5257\,
            in3 => \N__11887\,
            lcout => \U409_ADDRESS_DECODE.N_58_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.D_1_i_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8390\,
            in2 => \_gnd_net_\,
            in3 => \N__8868\,
            lcout => \D_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.CONFIGENn_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__7456\,
            in1 => \N__6533\,
            in2 => \N__5184\,
            in3 => \N__6624\,
            lcout => \CONFIGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.CONFIGENnC_net\,
            ce => 'H',
            sr => \N__11395\
        );

    \U409_AUTOCONFIG.LIDE_CONF_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__7449\,
            in1 => \N__6539\,
            in2 => \_gnd_net_\,
            in3 => \N__6617\,
            lcout => \U409_AUTOCONFIG.LIDE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__11394\
        );

    \U409_AUTOCONFIG.PRO_BASE_2_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5359\,
            in1 => \N__7906\,
            in2 => \N__8062\,
            in3 => \N__5166\,
            lcout => \PRO_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__11394\
        );

    \U409_AUTOCONFIG.PRO_BASE_0_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7904\,
            in1 => \N__5154\,
            in2 => \N__8152\,
            in3 => \N__5357\,
            lcout => \PRO_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__11394\
        );

    \U409_AUTOCONFIG.PRO_BASE_1_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__5358\,
            in1 => \N__7905\,
            in2 => \N__6754\,
            in3 => \N__5373\,
            lcout => \PRO_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_CONFC_net\,
            ce => 'H',
            sr => \N__11394\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_1_1_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5980\,
            in2 => \_gnd_net_\,
            in3 => \N__6849\,
            lcout => \U409_AUTOCONFIG.N_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_1_0_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5979\,
            in1 => \N__6215\,
            in2 => \N__6886\,
            in3 => \N__6112\,
            lcout => \U409_AUTOCONFIG.N_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIDEFO1_0_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__7467\,
            in1 => \N__8904\,
            in2 => \_gnd_net_\,
            in3 => \N__8778\,
            lcout => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1\,
            ltout => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7451\,
            in2 => \N__5362\,
            in3 => \N__6518\,
            lcout => \U409_AUTOCONFIG.CONFIGENn_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_0_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5347\,
            in1 => \N__6111\,
            in2 => \N__6885\,
            in3 => \N__6214\,
            lcout => \U409_AUTOCONFIG.N_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_A_14_2_0_a2_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__6213\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6110\,
            lcout => \U409_AUTOCONFIG.N_216_3\,
            ltout => \U409_AUTOCONFIG.N_216_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_o4_2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__5335\,
            in1 => \N__11875\,
            in2 => \N__5338\,
            in3 => \N__6912\,
            lcout => \U409_AUTOCONFIG.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_2_3_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__6997\,
            in1 => \N__7073\,
            in2 => \_gnd_net_\,
            in3 => \N__5670\,
            lcout => \U409_AUTOCONFIG.N_108\,
            ltout => \U409_AUTOCONFIG.N_108_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_3_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__6210\,
            in1 => \N__5737\,
            in2 => \N__5329\,
            in3 => \N__6045\,
            lcout => \U409_AUTOCONFIG.N_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.un1_AUTOVECTOR_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__5476\,
            in1 => \N__7123\,
            in2 => \N__5467\,
            in3 => \N__5449\,
            lcout => \U409_TRANSFER_ACK.un1_AUTOVECTOR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__5563\,
            in1 => \N__5443\,
            in2 => \N__5437\,
            in3 => \N__5578\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => \N__6279\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI9FMP_2_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7448\,
            in1 => \N__6337\,
            in2 => \_gnd_net_\,
            in3 => \N__5554\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_RNI9FMPZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIVV912_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__5788\,
            in1 => \N__6382\,
            in2 => \N__5425\,
            in3 => \N__7635\,
            lcout => \D_OUT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNISS912_1_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__6381\,
            in1 => \N__5569\,
            in2 => \N__7636\,
            in3 => \N__5524\,
            lcout => \D_OUT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_0_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010001"
        )
    port map (
            in0 => \N__5497\,
            in1 => \N__6307\,
            in2 => \N__5977\,
            in3 => \N__5617\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_0C_net\,
            ce => \N__6279\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_0_o2_2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__5962\,
            in1 => \N__6218\,
            in2 => \N__6118\,
            in3 => \N__5865\,
            lcout => \U409_AUTOCONFIG.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__6221\,
            in1 => \N__6116\,
            in2 => \_gnd_net_\,
            in3 => \N__5964\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__5386\,
            in1 => \N__6220\,
            in2 => \N__5380\,
            in3 => \N__5493\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.PR_OUT_1C_net\,
            ce => \N__6268\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_i_o4_0_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001100110011"
        )
    port map (
            in0 => \N__6219\,
            in1 => \N__11852\,
            in2 => \N__6887\,
            in3 => \N__5963\,
            lcout => \U409_AUTOCONFIG.N_91\,
            ltout => \U409_AUTOCONFIG.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001101"
        )
    port map (
            in0 => \N__6348\,
            in1 => \N__6850\,
            in2 => \N__5557\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.PR_OUT_1C_net\,
            ce => \N__6268\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000001010"
        )
    port map (
            in0 => \N__11853\,
            in1 => \N__5547\,
            in2 => \N__5629\,
            in3 => \N__5931\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => \N__6280\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_1_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000001100000"
        )
    port map (
            in0 => \N__5548\,
            in1 => \N__6928\,
            in2 => \N__5960\,
            in3 => \N__5613\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_7_i_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_1_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__11854\,
            in1 => \_gnd_net_\,
            in2 => \N__5539\,
            in3 => \_gnd_net_\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => \N__6280\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI7DMP_1_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__7455\,
            in1 => \N__5536\,
            in2 => \_gnd_net_\,
            in3 => \N__5530\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNI7DMPZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_3_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010101010"
        )
    port map (
            in0 => \N__11855\,
            in1 => \N__5515\,
            in2 => \N__6939\,
            in3 => \N__5935\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => \N__6280\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNO_0_2_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__6217\,
            in1 => \N__6932\,
            in2 => \N__5961\,
            in3 => \N__5492\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.PR_OUT_cnst_i_i_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_2_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001111"
        )
    port map (
            in0 => \N__5628\,
            in1 => \_gnd_net_\,
            in2 => \N__5791\,
            in3 => \N__6216\,
            lcout => \U409_AUTOCONFIG.PR_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_1C_net\,
            ce => \N__6280\,
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNIOGLSO_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__7099\,
            in1 => \N__6672\,
            in2 => \_gnd_net_\,
            in3 => \N__8421\,
            lcout => \PORTSIZE_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.un1_STATE_6_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__5675\,
            in1 => \N__6212\,
            in2 => \N__5755\,
            in3 => \N__6051\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_cnst_i_i_a2_0_3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7074\,
            in1 => \N__7003\,
            in2 => \N__5754\,
            in3 => \N__5674\,
            lcout => \U409_AUTOCONFIG.N_109\,
            ltout => \U409_AUTOCONFIG.N_109_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_cnst_i_i_a2_1_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6049\,
            in2 => \N__5632\,
            in3 => \N__6927\,
            lcout => \U409_AUTOCONFIG.N_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_i_a2_0_0_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6211\,
            in2 => \_gnd_net_\,
            in3 => \N__6050\,
            lcout => \U409_AUTOCONFIG.N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_2_0_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__5602\,
            in1 => \N__6142\,
            in2 => \N__6105\,
            in3 => \N__5939\,
            lcout => \U409_AUTOCONFIG.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_4_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__7516\,
            in1 => \N__9744\,
            in2 => \_gnd_net_\,
            in3 => \N__6496\,
            lcout => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_0_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10107\,
            in1 => \N__9913\,
            in2 => \N__10005\,
            in3 => \N__7798\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENnZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__8532\,
            in1 => \N__9729\,
            in2 => \N__5872\,
            in3 => \N__7734\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_2_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__7797\,
            in1 => \N__7733\,
            in2 => \N__6433\,
            in3 => \N__8101\,
            lcout => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_AUTOCONFIG_SPACE_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8867\,
            in2 => \_gnd_net_\,
            in3 => \N__8413\,
            lcout => \un1_AUTOCONFIG_SPACE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_3_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__11848\,
            in1 => \N__6934\,
            in2 => \N__5887\,
            in3 => \N__5869\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => \N__6278\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_3_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11849\,
            in2 => \_gnd_net_\,
            in3 => \N__5886\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_OUT_3C_net\,
            ce => \N__6278\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIH4AI_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7436\,
            lcout => \U409_AUTOCONFIG.D_OUT_sm0_0\,
            ltout => \U409_AUTOCONFIG.D_OUT_sm0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNI23A12_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__5803\,
            in1 => \N__5848\,
            in2 => \N__5839\,
            in3 => \N__7625\,
            lcout => \D_OUT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNIBHMP_3_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5815\,
            in1 => \N__5809\,
            in2 => \_gnd_net_\,
            in3 => \N__7438\,
            lcout => \U409_AUTOCONFIG.LIDE_OUT_RNIBHMPZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNI5BMP_0_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7437\,
            in1 => \N__5797\,
            in2 => \_gnd_net_\,
            in3 => \N__6286\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.LIDE_OUT_RNI5BMPZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.PR_OUT_RNIPP912_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__6391\,
            in1 => \N__7620\,
            in2 => \N__6385\,
            in3 => \N__6380\,
            lcout => \D_OUT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__7435\,
            in1 => \N__6534\,
            in2 => \N__6940\,
            in3 => \N__6955\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_2_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__6331\,
            in1 => \N__6349\,
            in2 => \N__6922\,
            in3 => \N__11850\,
            lcout => \U409_AUTOCONFIG.LIDE_OUTZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            ce => \N__6267\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_RNO_0_2_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6226\,
            in1 => \N__5978\,
            in2 => \N__6117\,
            in3 => \N__6894\,
            lcout => \U409_AUTOCONFIG.N_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_RNI04BC_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__6325\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6418\,
            lcout => \U409_AUTOCONFIG.STATE4\,
            ltout => \U409_AUTOCONFIG.STATE4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNI10V92_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111010101"
        )
    port map (
            in0 => \N__11851\,
            in1 => \N__6412\,
            in2 => \N__6310\,
            in3 => \N__8905\,
            lcout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_RNO_0_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000000"
        )
    port map (
            in0 => \N__6106\,
            in1 => \N__6225\,
            in2 => \N__6921\,
            in3 => \N__5968\,
            lcout => OPEN,
            ltout => \U409_AUTOCONFIG.N_103_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_OUT_0_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__6306\,
            in1 => \_gnd_net_\,
            in2 => \N__6289\,
            in3 => \N__11837\,
            lcout => \U409_AUTOCONFIG.BRIDGE_OUTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_OUT_2C_net\,
            ce => \N__6267\,
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_OUT_7_0_a2_3_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000000000"
        )
    port map (
            in0 => \N__6224\,
            in1 => \N__6084\,
            in2 => \N__6933\,
            in3 => \N__5950\,
            lcout => \U409_AUTOCONFIG.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_START_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__7624\,
            in1 => \N__10394\,
            in2 => \_gnd_net_\,
            in3 => \N__8417\,
            lcout => \U409_AUTOCONFIG.AC_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIJFAU_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8856\,
            in2 => \_gnd_net_\,
            in3 => \N__8782\,
            lcout => \U409_AUTOCONFIG.un1_PR_OUT_9_sqmuxa_0_a3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000010000"
        )
    port map (
            in0 => \N__7311\,
            in1 => \N__7360\,
            in2 => \N__11573\,
            in3 => \N__7285\,
            lcout => OPEN,
            ltout => \U409_CIA.CLK_CIA_r_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001101010"
        )
    port map (
            in0 => \N__11566\,
            in1 => \N__6466\,
            in2 => \N__6406\,
            in3 => \N__7338\,
            lcout => \CLK_CIA_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12844\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.un2_CIA_CLK_COUNT_cry_1_c_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7251\,
            in2 => \N__7228\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_12_0_\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_2_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7359\,
            in2 => \_gnd_net_\,
            in3 => \N__6403\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_2\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_1\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7260\,
            in1 => \N__7306\,
            in2 => \_gnd_net_\,
            in3 => \N__6400\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_3\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_2\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_4_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7284\,
            in2 => \_gnd_net_\,
            in3 => \N__6397\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_4\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_3\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_5_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__7261\,
            in1 => \N__7336\,
            in2 => \_gnd_net_\,
            in3 => \N__6394\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_5\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_4\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_6_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7174\,
            in2 => \_gnd_net_\,
            in3 => \N__6472\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_6\,
            ltout => OPEN,
            carryin => \U409_CIA.un2_CIA_CLK_COUNT_cry_5\,
            carryout => \U409_CIA.un2_CIA_CLK_COUNT_cry_6\,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_7_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7191\,
            in2 => \_gnd_net_\,
            in3 => \N__6469\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12846\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CLK_CIA_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__7252\,
            in1 => \N__7173\,
            in2 => \N__7192\,
            in3 => \N__7224\,
            lcout => \U409_CIA.CLK_CIA6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_3_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__10016\,
            in1 => \N__10108\,
            in2 => \N__7993\,
            in3 => \N__6487\,
            lcout => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RTC_ENn_i_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__8543\,
            in1 => \N__6460\,
            in2 => \N__9760\,
            in3 => \N__7723\,
            lcout => \U409_ADDRESS_DECODE_un1_RTC_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_BASE_1_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__7874\,
            in1 => \N__7493\,
            in2 => \N__8137\,
            in3 => \N__7747\,
            lcout => \LIDE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_2_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7873\,
            in1 => \N__6429\,
            in2 => \N__6752\,
            in3 => \N__8014\,
            lcout => \BRIDGE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.LIDE_BASE_2_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__7494\,
            in1 => \N__7875\,
            in2 => \N__7657\,
            in3 => \N__6744\,
            lcout => \LIDE_BASE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.LIDE_BASE_5_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7971\,
            in1 => \N__7876\,
            in2 => \N__8138\,
            in3 => \N__7549\,
            lcout => \LIDE_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.LIDE_BASE_6_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__7877\,
            in1 => \N__7972\,
            in2 => \N__7564\,
            in3 => \N__6745\,
            lcout => \LIDE_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.CONFIGURED_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__6544\,
            in1 => \N__6628\,
            in2 => \N__7450\,
            in3 => \N__7612\,
            lcout => \CONFIGURED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.LIDE_BASE_1C_net\,
            ce => 'H',
            sr => \N__11393\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_0_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7865\,
            in1 => \N__6600\,
            in2 => \N__7953\,
            in3 => \N__8011\,
            lcout => \BRIDGE_BASE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_0C_net\,
            ce => 'H',
            sr => \N__11392\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__6923\,
            in1 => \N__7406\,
            in2 => \_gnd_net_\,
            in3 => \N__6953\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FUZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000001000"
        )
    port map (
            in0 => \N__7613\,
            in1 => \N__9395\,
            in2 => \N__9301\,
            in3 => \N__6601\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_i_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__6592\,
            in1 => \N__6583\,
            in2 => \N__6574\,
            in3 => \N__6571\,
            lcout => \U409_ADDRESS_DECODE_un1_BREG_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2_1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7407\,
            in1 => \N__6543\,
            in2 => \N__6938\,
            in3 => \N__6954\,
            lcout => \U409_AUTOCONFIG.LIDE_CONF_RNIUIPA2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_BREG_ENn_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010000100001"
        )
    port map (
            in0 => \N__9899\,
            in1 => \N__10209\,
            in2 => \N__6688\,
            in3 => \N__7084\,
            lcout => \U409_ADDRESS_DECODE.un1_BREG_ENnZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_4_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__7888\,
            in1 => \N__6483\,
            in2 => \N__7954\,
            in3 => \N__7529\,
            lcout => \BRIDGE_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net\,
            ce => 'H',
            sr => \N__11388\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_7_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7530\,
            in1 => \N__7890\,
            in2 => \N__8061\,
            in3 => \N__7083\,
            lcout => \BRIDGE_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net\,
            ce => 'H',
            sr => \N__11388\
        );

    \U409_AUTOCONFIG.STATE_RNIU6QK1_0_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7075\,
            in1 => \N__7018\,
            in2 => \N__6970\,
            in3 => \N__8920\,
            lcout => \U409_AUTOCONFIG.un1_STATE_6_0\,
            ltout => \U409_AUTOCONFIG.un1_STATE_6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1_0_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__6864\,
            in1 => \_gnd_net_\,
            in2 => \N__6757\,
            in3 => \N__7427\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0\,
            ltout => \U409_AUTOCONFIG.BRIDGE_CONF_RNID7FU1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_6_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__7889\,
            in1 => \N__6753\,
            in2 => \N__6691\,
            in3 => \N__6684\,
            lcout => \BRIDGE_BASE_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_4C_net\,
            ce => 'H',
            sr => \N__11388\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8205\,
            in2 => \_gnd_net_\,
            in3 => \N__8191\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__8673\
        );

    \U409_CIA.VMA_RNO_0_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__7366\,
            in1 => \N__7337\,
            in2 => \N__7312\,
            in3 => \N__7159\,
            lcout => OPEN,
            ltout => \U409_CIA.VMA_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__6676\,
            in1 => \N__10904\,
            in2 => \N__6658\,
            in3 => \N__7225\,
            lcout => \U409_CIA.VMAZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_0_0_0_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__9895\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10090\,
            lcout => \U409_ADDRESS_DECODE.un1_RTC_ENn_2\,
            ltout => \U409_ADDRESS_DECODE.un1_RTC_ENn_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_i_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__8496\,
            in1 => \N__8544\,
            in2 => \N__6655\,
            in3 => \N__9708\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNO_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000101000"
        )
    port map (
            in0 => \N__7248\,
            in1 => \N__7282\,
            in2 => \N__7226\,
            in3 => \N__7358\,
            lcout => \U409_CIA.un1_CIA_CLK_COUNT_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIGOMD1_2_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7357\,
            in1 => \N__7214\,
            in2 => \N__7339\,
            in3 => \N__7247\,
            lcout => OPEN,
            ltout => \U409_CIA.CIA_CLK_COUNT11_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNICTDR2_3_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__7307\,
            in1 => \N__7283\,
            in2 => \N__7264\,
            in3 => \N__7158\,
            lcout => \U409_CIA.CIA_CLK_COUNT11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_0_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7249\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__7250\,
            in1 => \_gnd_net_\,
            in2 => \N__7227\,
            in3 => \_gnd_net_\,
            lcout => \U409_CIA.CIA_CLK_COUNTZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12845\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.CIA_CLK_COUNT_RNIHLRM_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7187\,
            in2 => \_gnd_net_\,
            in3 => \N__7172\,
            lcout => \U409_CIA.CLK_CIA6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m20_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9398\,
            in1 => \N__9758\,
            in2 => \N__9100\,
            in3 => \N__10017\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.N_77_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_22_0_i_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10111\,
            in2 => \N__7147\,
            in3 => \_gnd_net_\,
            lcout => \N_22_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNIO8F0F_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__7116\,
            in1 => \N__8357\,
            in2 => \N__8743\,
            in3 => \N__8343\,
            lcout => \U409_ADDRESS_DECODE.PORTSIZE_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_0_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001001000001"
        )
    port map (
            in0 => \N__7813\,
            in1 => \N__7746\,
            in2 => \N__7732\,
            in3 => \N__7653\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7570\,
            in1 => \N__7537\,
            in2 => \N__7642\,
            in3 => \N__8428\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0\,
            ltout => \U409_ADDRESS_DECODE.ATA_SPACEZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000100000"
        )
    port map (
            in0 => \N__11815\,
            in1 => \N__8866\,
            in2 => \N__7639\,
            in3 => \N__8342\,
            lcout => \U409_ADDRESS_DECODE.ATA_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__11175\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_3_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__9396\,
            in1 => \N__10214\,
            in2 => \N__8080\,
            in3 => \N__7608\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__9914\,
            in1 => \N__7560\,
            in2 => \N__9754\,
            in3 => \N__7548\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_5_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__8148\,
            in1 => \N__7909\,
            in2 => \N__7512\,
            in3 => \N__7531\,
            lcout => \BRIDGE_BASE_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.LIDE_BASE_3_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__7910\,
            in1 => \N__7495\,
            in2 => \N__8443\,
            in3 => \N__8047\,
            lcout => \LIDE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.BRIDGE_CONF_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__7477\,
            in1 => \N__7428\,
            in2 => \_gnd_net_\,
            in3 => \N__8919\,
            lcout => \U409_AUTOCONFIG.BRIDGE_CONFZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_1_LC_10_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__8147\,
            in1 => \N__8012\,
            in2 => \N__8097\,
            in3 => \N__7907\,
            lcout => \BRIDGE_BASE_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.LIDE_BASE_7_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7970\,
            in1 => \N__8048\,
            in2 => \N__7918\,
            in3 => \N__8076\,
            lcout => \LIDE_BASE_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.BRIDGE_BASE_3_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__8046\,
            in1 => \N__8013\,
            in2 => \N__7989\,
            in3 => \N__7908\,
            lcout => \BRIDGE_BASE_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_AUTOCONFIG.LIDE_BASE_4_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__7969\,
            in1 => \N__7952\,
            in2 => \N__7917\,
            in3 => \N__8455\,
            lcout => \LIDE_BASE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.BRIDGE_BASE_5C_net\,
            ce => 'H',
            sr => \N__11389\
        );

    \U409_ADDRESS_DECODE.m33_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8242\,
            in1 => \N__8565\,
            in2 => \N__8311\,
            in3 => \N__7819\,
            lcout => \N_71_mux\,
            ltout => \N_71_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m38_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001110100111111"
        )
    port map (
            in0 => \N__11498\,
            in1 => \N__8976\,
            in2 => \N__7825\,
            in3 => \N__8942\,
            lcout => \N_23\,
            ltout => \N_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8223\,
            in2 => \N__7822\,
            in3 => \N__8567\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8674\
        );

    \U409_ADDRESS_DECODE.m33_3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8221\,
            in1 => \N__8187\,
            in2 => \N__8595\,
            in3 => \N__8269\,
            lcout => \U409_ADDRESS_DECODE.m33Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m27_3_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8188\,
            in1 => \N__8222\,
            in2 => \N__8275\,
            in3 => \N__8586\,
            lcout => OPEN,
            ltout => \U409_ADDRESS_DECODE.m27Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m27_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__8566\,
            in1 => \N__8308\,
            in2 => \N__8287\,
            in3 => \N__8243\,
            lcout => \N_70_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_7_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000010000000"
        )
    port map (
            in0 => \N__8284\,
            in1 => \N__8979\,
            in2 => \N__8623\,
            in3 => \N__8309\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8674\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_6_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__8978\,
            in1 => \N__8283\,
            in2 => \_gnd_net_\,
            in3 => \N__8619\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_1C_net\,
            ce => 'H',
            sr => \N__8674\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI11UH2_5_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__8244\,
            in1 => \N__8254\,
            in2 => \N__8206\,
            in3 => \N__8190\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__8274\,
            in1 => \N__8160\,
            in2 => \N__8596\,
            in3 => \N__8621\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__8656\
        );

    \U409_ADDRESS_DECODE.m33_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8590\,
            in2 => \_gnd_net_\,
            in3 => \N__8273\,
            lcout => \U409_ADDRESS_DECODE_m33_1\,
            ltout => \U409_ADDRESS_DECODE_m33_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_5_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110101000000000"
        )
    port map (
            in0 => \N__8245\,
            in1 => \N__8161\,
            in2 => \N__8248\,
            in3 => \N__8622\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__8656\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNI7S9R_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8568\,
            in2 => \_gnd_net_\,
            in3 => \N__8224\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_RNISRU81_2_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8189\,
            in2 => \N__8164\,
            in3 => \_gnd_net_\,
            lcout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3\,
            ltout => \U409_TRANSFER_ACK.un1_DELAYED_TACK_COUNTER_2_c3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_3_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__8620\,
            in1 => \_gnd_net_\,
            in2 => \N__8599\,
            in3 => \N__8591\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__8656\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER_0_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011001010101"
        )
    port map (
            in0 => \N__8569\,
            in1 => \N__8980\,
            in2 => \N__11497\,
            in3 => \N__8944\,
            lcout => \U409_TRANSFER_ACK_DELAYED_TACK_COUNTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_COUNTER_4C_net\,
            ce => 'H',
            sr => \N__8656\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_COUNTER16_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10395\,
            in2 => \_gnd_net_\,
            in3 => \N__11202\,
            lcout => \N_52_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_REGSPACEn_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10245\,
            in1 => \N__8548\,
            in2 => \N__8503\,
            in3 => \N__9724\,
            lcout => \U409_ADDRESS_DECODE_un1_REGSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_SPACE_1_0_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000000001001"
        )
    port map (
            in0 => \N__10110\,
            in1 => \N__8454\,
            in2 => \N__10009\,
            in3 => \N__8439\,
            lcout => \U409_ADDRESS_DECODE.ATA_SPACE_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.LV_SPACE_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__8742\,
            in1 => \N__8688\,
            in2 => \N__8362\,
            in3 => \N__8422\,
            lcout => \BUFENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ATA_EN_RNITH4D5_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8358\,
            in2 => \_gnd_net_\,
            in3 => \N__8344\,
            lcout => \U409_ADDRESS_DECODE_un1_ATA_ENn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8310\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.DELAYED_TACK_EN_nerC_net\,
            ce => \N__8926\,
            sr => \N__8666\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__9018\,
            in1 => \N__9399\,
            in2 => \N__10219\,
            in3 => \N__9796\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_1_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000011000000"
        )
    port map (
            in0 => \N__8837\,
            in1 => \N__8895\,
            in2 => \N__11836\,
            in3 => \N__8770\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_0_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__8769\,
            in1 => \N__11788\,
            in2 => \N__8903\,
            in3 => \N__8989\,
            lcout => \U409_AUTOCONFIG.STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.STATE_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_sbtinv_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8977\,
            in2 => \N__8953\,
            in3 => \N__8943\,
            lcout => \U409_TRANSFER_ACK.N_20_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.STATE_RNIF4QU_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8891\,
            in2 => \_gnd_net_\,
            in3 => \N__8768\,
            lcout => \U409_AUTOCONFIG.STATE_d_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_AUTOCONFIG.AC_TACK_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111010001000"
        )
    port map (
            in0 => \N__9522\,
            in1 => \N__8902\,
            in2 => \N__8869\,
            in3 => \N__8777\,
            lcout => \AC_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_AUTOCONFIG.AC_TACKC_net\,
            ce => 'H',
            sr => \N__11383\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_i_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__8726\,
            in1 => \N__8710\,
            in2 => \N__8692\,
            in3 => \N__11795\,
            lcout => \U409_TRANSFER_ACK.DELAYED_TACK_RST_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_1_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9912\,
            in2 => \_gnd_net_\,
            in3 => \N__9723\,
            lcout => \U409_ADDRESS_DECODE.N_60_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_CLK40_IN_c_g_THRU_LUT4_0_LC_12_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11206\,
            lcout => \GB_BUFFER_CLK40_IN_c_g_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS0_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9296\,
            in1 => \N__9237\,
            in2 => \N__9215\,
            in3 => \N__9150\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.CS1_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9297\,
            in1 => \N__9238\,
            in2 => \N__9216\,
            in3 => \N__9151\,
            lcout => \U409_ADDRESS_DECODE.CSZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS1n_i_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__9217\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9160\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS1n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_CIA.VMA_RNI692L_0_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11731\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10924\,
            lcout => \CIA_ENABLE\,
            ltout => \CIA_ENABLE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_CIACS0n_i_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9154\,
            in3 => \N__9141\,
            lcout => \U409_ADDRESS_DECODE_un1_CIACS0n_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.N_77_mux_i_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__9403\,
            in1 => \N__9096\,
            in2 => \N__10010\,
            in3 => \N__9759\,
            lcout => \N_77_mux_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.un1_RAMSPACEn_i_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011111"
        )
    port map (
            in0 => \N__9397\,
            in1 => \N__9785\,
            in2 => \N__9025\,
            in3 => \N__10190\,
            lcout => \U409_ADDRESS_DECODE_un1_RAMSPACEn_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_0_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__9450\,
            in1 => \N__9432\,
            in2 => \N__11775\,
            in3 => \N__9414\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_COUNTER_1_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__9431\,
            in1 => \N__11738\,
            in2 => \_gnd_net_\,
            in3 => \N__9449\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.DELAYED_TACK_EN_ner_RNIKDE9_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9529\,
            in2 => \_gnd_net_\,
            in3 => \N__10332\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER5_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_RNIFT8M_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__9523\,
            in1 => \N__10939\,
            in2 => \N__9508\,
            in3 => \N__10314\,
            lcout => \U409_TRANSFER_ACK.TACK_COUNTER6\,
            ltout => \U409_TRANSFER_ACK.TACK_COUNTER6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_RNO_0_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000111011101"
        )
    port map (
            in0 => \N__9448\,
            in1 => \N__9430\,
            in2 => \N__9505\,
            in3 => \N__9469\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.TACK_OUTn_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_OUTn_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__9470\,
            in1 => \_gnd_net_\,
            in2 => \N__9502\,
            in3 => \N__11739\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010011001"
        )
    port map (
            in0 => \N__10888\,
            in1 => \N__10806\,
            in2 => \_gnd_net_\,
            in3 => \N__11463\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__11382\
        );

    \U409_TRANSFER_ACK.TACK_EN_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000001110001"
        )
    port map (
            in0 => \N__9451\,
            in1 => \N__9433\,
            in2 => \N__9589\,
            in3 => \N__9415\,
            lcout => \TACK_EN\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__11382\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011000000"
        )
    port map (
            in0 => \N__10024\,
            in1 => \N__9388\,
            in2 => \N__10234\,
            in3 => \N__9622\,
            lcout => \ROMEN\,
            ltout => \ROMEN_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIRHPR5_0_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9307\,
            in3 => \N__11434\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_RNO_0_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10755\,
            in1 => \N__10805\,
            in2 => \N__9304\,
            in3 => \N__10858\,
            lcout => \U409_TRANSFER_ACK.un1_ROM_TACK_COUNTER20_3_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_0_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9740\,
            in1 => \N__10252\,
            in2 => \N__10218\,
            in3 => \N__10011\,
            lcout => \U409_ADDRESS_DECODE.N_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIV1RD_3_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010111011"
        )
    port map (
            in0 => \N__10647\,
            in1 => \N__10715\,
            in2 => \_gnd_net_\,
            in3 => \N__10754\,
            lcout => \U409_TRANSFER_ACK.N_42_i\,
            ltout => \U409_TRANSFER_ACK.N_42_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_2_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000001100000"
        )
    port map (
            in0 => \N__11435\,
            in1 => \N__10648\,
            in2 => \N__10222\,
            in3 => \N__10707\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_1_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__10213\,
            in1 => \N__10109\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.ROMEN_0_a3_2_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__10012\,
            in1 => \N__9916\,
            in2 => \N__9795\,
            in3 => \N__9728\,
            lcout => \U409_ADDRESS_DECODE.ROMEN_0_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.TACK_EN_RNIPUKQ5_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9616\,
            in2 => \_gnd_net_\,
            in3 => \N__9590\,
            lcout => \TCIn_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11796\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_LC_13_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__10425\,
            in1 => \N__11203\,
            in2 => \N__10407\,
            in3 => \N__10348\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTERZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__11386\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_RNO_0_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__10426\,
            in1 => \_gnd_net_\,
            in2 => \N__10408\,
            in3 => \N__11842\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.IRQ_TACK_COUNTER_0_sqmuxa_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.IRQ_TACK_EN_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__11204\,
            in1 => \N__10347\,
            in2 => \N__10336\,
            in3 => \N__10333\,
            lcout => \U409_TRANSFER_ACK.IRQ_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.IRQ_TACK_COUNTERC_net\,
            ce => 'H',
            sr => \N__11386\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__10321\,
            in1 => \N__10315\,
            in2 => \N__10726\,
            in3 => \N__10258\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11385\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_3_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100000010"
        )
    port map (
            in0 => \N__10807\,
            in1 => \N__11459\,
            in2 => \N__10887\,
            in3 => \N__10759\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11385\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_1_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__11458\,
            in1 => \N__10859\,
            in2 => \_gnd_net_\,
            in3 => \N__11440\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11385\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNI87LI_2_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000010"
        )
    port map (
            in0 => \N__10646\,
            in1 => \N__10795\,
            in2 => \N__10717\,
            in3 => \N__10848\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_NE_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIGEA51_3_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000010000"
        )
    port map (
            in0 => \N__10602\,
            in1 => \N__11436\,
            in2 => \N__10303\,
            in3 => \N__10756\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0\,
            ltout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER23_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROMENn_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111010011111100"
        )
    port map (
            in0 => \N__11505\,
            in1 => \N__10275\,
            in2 => \N__10300\,
            in3 => \N__10297\,
            lcout => \ROMENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROMENnC_net\,
            ce => 'H',
            sr => \N__11384\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_0_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__10861\,
            in1 => \N__10867\,
            in2 => \N__10808\,
            in3 => \N__10264\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m43_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__10489\,
            in1 => \N__10510\,
            in2 => \_gnd_net_\,
            in3 => \N__10534\,
            lcout => \PCIAT_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.m45_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__10533\,
            in1 => \N__10509\,
            in2 => \_gnd_net_\,
            in3 => \N__10482\,
            lcout => \PCIAT_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un3_COUNTER60_1_cry_1_c_LC_14_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11315\,
            in2 => \N__10963\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_6_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_2_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11334\,
            in2 => \_gnd_net_\,
            in3 => \N__10444\,
            lcout => \U409_TICK.COUNTER60Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_1\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_2\,
            clk => \N__12598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_3_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11265\,
            in2 => \_gnd_net_\,
            in3 => \N__10441\,
            lcout => \U409_TICK.COUNTER60Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_2\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_3\,
            clk => \N__12598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_4_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11067\,
            in2 => \_gnd_net_\,
            in3 => \N__10438\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_3\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_5_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11085\,
            in2 => \_gnd_net_\,
            in3 => \N__10435\,
            lcout => \U409_TICK.COUNTER60Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_4\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_5\,
            clk => \N__12598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_6_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11016\,
            in2 => \_gnd_net_\,
            in3 => \N__10432\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_5\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_7_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10977\,
            in2 => \_gnd_net_\,
            in3 => \N__10429\,
            lcout => \U409_TICK.COUNTER60Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_6\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_7\,
            clk => \N__12598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_8_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__11044\,
            in3 => \N__10582\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_7\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_9_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11055\,
            in2 => \_gnd_net_\,
            in3 => \N__10579\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_14_7_0_\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_10_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10992\,
            in2 => \_gnd_net_\,
            in3 => \N__10576\,
            lcout => \U409_TICK.COUNTER60Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_9\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_10\,
            clk => \N__12599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_11_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11280\,
            in2 => \_gnd_net_\,
            in3 => \N__10573\,
            lcout => \U409_TICK.COUNTER60Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_10\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_11\,
            clk => \N__12599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_12_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11346\,
            in2 => \_gnd_net_\,
            in3 => \N__10570\,
            lcout => \U409_TICK.COUNTER60Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_11\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_12\,
            clk => \N__12599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_13_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11004\,
            in2 => \_gnd_net_\,
            in3 => \N__10567\,
            lcout => \U409_TICK.COUNTER60Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_12\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_13\,
            clk => \N__12599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_14_LC_14_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11244\,
            in2 => \_gnd_net_\,
            in3 => \N__10564\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_13\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNO_0_15_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11220\,
            in2 => \_gnd_net_\,
            in3 => \N__10561\,
            lcout => \U409_TICK.COUNTER60_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un3_COUNTER60_1_cry_14\,
            carryout => \U409_TICK.un3_COUNTER60_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_16_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11299\,
            in2 => \_gnd_net_\,
            in3 => \N__10558\,
            lcout => \U409_TICK.COUNTER60Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12599\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_TACK_EN_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001001100"
        )
    port map (
            in0 => \N__11627\,
            in1 => \N__10938\,
            in2 => \N__11650\,
            in3 => \N__11116\,
            lcout => \U409_TRANSFER_ACK.CIA_TACK_ENZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11390\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_1_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11911\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11390\
        );

    \U409_TRANSFER_ACK.CIA_ENABLED_0_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10923\,
            lcout => \U409_TRANSFER_ACK.CIA_ENABLEDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_TACK_ENC_net\,
            ce => 'H',
            sr => \N__11390\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNO_0_0_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010100"
        )
    port map (
            in0 => \N__11430\,
            in1 => \N__10812\,
            in2 => \N__10860\,
            in3 => \N__10758\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER_6_f0_0_a2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_RNIJBK9_0_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10851\,
            in2 => \_gnd_net_\,
            in3 => \N__11429\,
            lcout => \U409_TRANSFER_ACK.N_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_3_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100001010000100"
        )
    port map (
            in0 => \N__10637\,
            in1 => \N__10849\,
            in2 => \N__10716\,
            in3 => \N__11420\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_NE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_EN_RNO_1_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000110000010"
        )
    port map (
            in0 => \N__10850\,
            in1 => \N__10813\,
            in2 => \N__10603\,
            in3 => \N__10757\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTER22_NE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER21_0_i_0_x3_0_0_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10708\,
            in2 => \_gnd_net_\,
            in3 => \N__10628\,
            lcout => \U409_TRANSFER_ACK.N_31_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_9_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12049\,
            in1 => \N__12122\,
            in2 => \N__12090\,
            in3 => \N__10588\,
            lcout => \U409_TICK.COUNTER60Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_8_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__12121\,
            in1 => \N__12051\,
            in2 => \N__11095\,
            in3 => \N__12086\,
            lcout => \U409_TICK.COUNTER60Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_1_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10961\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11319\,
            lcout => \U409_TICK.COUNTER60Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIHJU51_4_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__11086\,
            in1 => \N__10960\,
            in2 => \_gnd_net_\,
            in3 => \N__11068\,
            lcout => \U409_TICK.TICK603_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_4_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__11074\,
            in1 => \N__12082\,
            in2 => \N__12124\,
            in3 => \N__12052\,
            lcout => \U409_TICK.COUNTER60Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNICDC71_14_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11056\,
            in1 => \N__11043\,
            in2 => \N__11020\,
            in3 => \N__11245\,
            lcout => \U409_TICK.TICK603_9\,
            ltout => \U409_TICK.TICK603_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_6_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12120\,
            in1 => \N__12050\,
            in2 => \N__11029\,
            in3 => \N__11026\,
            lcout => \U409_TICK.COUNTER60Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12600\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI2USG_10_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__11005\,
            in1 => \N__10993\,
            in2 => \N__10981\,
            in3 => \N__11221\,
            lcout => \U409_TICK.TICK603_10\,
            ltout => \U409_TICK.TICK603_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_0_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001111111"
        )
    port map (
            in0 => \N__12079\,
            in1 => \N__12053\,
            in2 => \N__10966\,
            in3 => \N__10962\,
            lcout => \U409_TICK.COUNTER60Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNIDB4S_16_LC_15_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11347\,
            in1 => \N__11335\,
            in2 => \N__11323\,
            in3 => \N__11298\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK603_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_RNI335G2_11_LC_15_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11287\,
            in1 => \N__11281\,
            in2 => \N__11269\,
            in3 => \N__11266\,
            lcout => \U409_TICK.TICK603_14\,
            ltout => \U409_TICK.TICK603_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_14_LC_15_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12115\,
            in1 => \N__12081\,
            in2 => \N__11254\,
            in3 => \N__11251\,
            lcout => \U409_TICK.COUNTER60Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER60_15_LC_15_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__12080\,
            in1 => \N__12116\,
            in2 => \N__11233\,
            in3 => \N__12054\,
            lcout => \U409_TICK.COUNTER60Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_0_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011111110111"
        )
    port map (
            in0 => \N__11921\,
            in1 => \N__11909\,
            in2 => \N__11628\,
            in3 => \N__11115\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.CIA_STATE_RNO_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_0_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001010001010"
        )
    port map (
            in0 => \N__11846\,
            in1 => \N__11649\,
            in2 => \N__11209\,
            in3 => \N__11101\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNI9HNJ_1_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11541\,
            in1 => \N__11601\,
            in2 => \_gnd_net_\,
            in3 => \N__11205\,
            lcout => \U409_TRANSFER_ACK.N_17_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_RNIHJ5G_1_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11540\,
            lcout => \U409_TRANSFER_ACK.N_3_0\,
            ltout => \U409_TRANSFER_ACK.N_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_1_0_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__11908\,
            in1 => \N__11625\,
            in2 => \N__11104\,
            in3 => \N__11923\,
            lcout => \U409_TRANSFER_ACK.CIA_STATE_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_RNO_0_1_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000011111"
        )
    port map (
            in0 => \N__11922\,
            in1 => \N__11910\,
            in2 => \N__11629\,
            in3 => \N__11893\,
            lcout => OPEN,
            ltout => \U409_TRANSFER_ACK.N_55_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.CIA_STATE_1_LC_15_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101000001000"
        )
    port map (
            in0 => \N__11847\,
            in1 => \N__11648\,
            in2 => \N__11632\,
            in3 => \N__11626\,
            lcout => \U409_TRANSFER_ACK.CIA_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.CIA_STATE_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TRANSFER_ACK.LASTCLK_1_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11542\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__11391\
        );

    \U409_TRANSFER_ACK.LASTCLK_0_LC_15_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11586\,
            lcout => \U409_TRANSFER_ACK.LASTCLKZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.LASTCLK_1C_net\,
            ce => 'H',
            sr => \N__11391\
        );

    \U409_TRANSFER_ACK.ROM_TACK_COUNTER_0_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__11527\,
            in1 => \N__11518\,
            in2 => \N__11512\,
            in3 => \N__11464\,
            lcout => \U409_TRANSFER_ACK.ROM_TACK_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU409_TRANSFER_ACK.ROM_TACK_COUNTER_0C_net\,
            ce => 'H',
            sr => \N__11387\
        );

    \U409_TICK.COUNTER50_15_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111000011110000"
        )
    port map (
            in0 => \N__12733\,
            in1 => \N__12704\,
            in2 => \N__12775\,
            in3 => \N__12660\,
            lcout => \U409_TICK.COUNTER50Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_13_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12702\,
            in1 => \N__12734\,
            in2 => \N__12668\,
            in3 => \N__12286\,
            lcout => \U409_TICK.COUNTER50Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_9_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12705\,
            in1 => \N__12736\,
            in2 => \N__12669\,
            in3 => \N__12346\,
            lcout => \U409_TICK.COUNTER50Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNII24V_14_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__12388\,
            in1 => \N__12811\,
            in2 => \N__12166\,
            in3 => \N__12787\,
            lcout => \U409_TICK.TICK503_10\,
            ltout => \U409_TICK.TICK503_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_14_LC_16_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12703\,
            in1 => \N__12735\,
            in2 => \N__12127\,
            in3 => \N__12796\,
            lcout => \U409_TICK.COUNTER50Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12601\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK60_LC_16_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12123\,
            in1 => \N__12012\,
            in2 => \N__12091\,
            in3 => \N__12055\,
            lcout => \TICK60_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_1_LC_16_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__12226\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12246\,
            lcout => \U409_TICK.COUNTER50Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12604\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_17_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNID6CP_3_LC_17_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__12148\,
            in1 => \N__12181\,
            in2 => \_gnd_net_\,
            in3 => \N__12220\,
            lcout => \U409_TICK.TICK503_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIUHF01_16_LC_17_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12373\,
            in1 => \N__12247\,
            in2 => \N__12199\,
            in3 => \N__12757\,
            lcout => OPEN,
            ltout => \U409_TICK.TICK503_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNITU182_10_LC_17_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__11935\,
            in1 => \N__12316\,
            in2 => \N__11929\,
            in3 => \N__12337\,
            lcout => \U409_TICK.TICK503_14\,
            ltout => \U409_TICK.TICK503_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_6_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010101010101010"
        )
    port map (
            in0 => \N__12397\,
            in1 => \N__12697\,
            in2 => \N__11926\,
            in3 => \N__12663\,
            lcout => \U409_TICK.COUNTER50Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.TICK50_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__12661\,
            in1 => \N__12738\,
            in2 => \N__12706\,
            in3 => \N__12261\,
            lcout => \TICK50_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_0_LC_17_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__12221\,
            in1 => \N__12696\,
            in2 => \N__12742\,
            in3 => \N__12662\,
            lcout => \U409_TICK.COUNTER50Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNIH14V_11_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__12298\,
            in1 => \N__12358\,
            in2 => \N__12415\,
            in3 => \N__12619\,
            lcout => \U409_TICK.TICK503_9\,
            ltout => \U409_TICK.TICK503_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_5_LC_17_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__12737\,
            in1 => \N__12136\,
            in2 => \N__12250\,
            in3 => \N__12664\,
            lcout => \U409_TICK.COUNTER50Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12602\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.un2_COUNTER50_1_cry_1_c_LC_17_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12242\,
            in2 => \N__12225\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_17_5_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_2_LC_17_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12195\,
            in2 => \_gnd_net_\,
            in3 => \N__12184\,
            lcout => \U409_TICK.COUNTER50Z0Z_2\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_1\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_2\,
            clk => \N__12605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_3_LC_17_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12180\,
            in2 => \_gnd_net_\,
            in3 => \N__12169\,
            lcout => \U409_TICK.COUNTER50Z0Z_3\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_2\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_3\,
            clk => \N__12605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_4_LC_17_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12162\,
            in2 => \_gnd_net_\,
            in3 => \N__12151\,
            lcout => \U409_TICK.COUNTER50Z0Z_4\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_3\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_4\,
            clk => \N__12605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_5_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12147\,
            in2 => \_gnd_net_\,
            in3 => \N__12130\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_4\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_6_LC_17_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12414\,
            in3 => \N__12391\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_5\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_7_LC_17_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12387\,
            in2 => \_gnd_net_\,
            in3 => \N__12376\,
            lcout => \U409_TICK.COUNTER50Z0Z_7\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_6\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_7\,
            clk => \N__12605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_8_LC_17_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12372\,
            in2 => \_gnd_net_\,
            in3 => \N__12361\,
            lcout => \U409_TICK.COUNTER50Z0Z_8\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_7\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_8\,
            clk => \N__12605\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_9_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12357\,
            in2 => \_gnd_net_\,
            in3 => \N__12340\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_9\,
            ltout => OPEN,
            carryin => \bfn_17_6_0_\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_10_LC_17_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12333\,
            in2 => \_gnd_net_\,
            in3 => \N__12322\,
            lcout => \U409_TICK.COUNTER50Z0Z_10\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_9\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_10\,
            clk => \N__12606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_11_LC_17_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12618\,
            in2 => \_gnd_net_\,
            in3 => \N__12319\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_11\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_10\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_12_LC_17_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12312\,
            in2 => \_gnd_net_\,
            in3 => \N__12301\,
            lcout => \U409_TICK.COUNTER50Z0Z_12\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_11\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_12\,
            clk => \N__12606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_13_LC_17_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12297\,
            in2 => \_gnd_net_\,
            in3 => \N__12280\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_13\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_12\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_14_LC_17_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12810\,
            in2 => \_gnd_net_\,
            in3 => \N__12790\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_14\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_13\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_RNO_0_15_LC_17_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12786\,
            in2 => \_gnd_net_\,
            in3 => \N__12763\,
            lcout => \U409_TICK.COUNTER50_RNO_0Z0Z_15\,
            ltout => OPEN,
            carryin => \U409_TICK.un2_COUNTER50_1_cry_14\,
            carryout => \U409_TICK.un2_COUNTER50_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_16_LC_17_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12756\,
            in2 => \_gnd_net_\,
            in3 => \N__12760\,
            lcout => \U409_TICK.COUNTER50Z0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12606\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_TICK.COUNTER50_11_LC_18_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111100000000"
        )
    port map (
            in0 => \N__12732\,
            in1 => \N__12701\,
            in2 => \N__12670\,
            in3 => \N__12625\,
            lcout => \U409_TICK.COUNTER50Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__12607\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS0_LC_19_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12471\,
            lcout => \PCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS1_LC_19_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__12472\,
            in1 => \N__12486\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \SCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.PCS1_LC_20_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12532\,
            in2 => \_gnd_net_\,
            in3 => \N__12469\,
            lcout => \PCS1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U409_ADDRESS_DECODE.SCS0_LC_20_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12487\,
            in2 => \_gnd_net_\,
            in3 => \N__12470\,
            lcout => \SCS0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AGNUS_CLK_obuf_RNO_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12874\,
            in1 => \N__12862\,
            in2 => \_gnd_net_\,
            in3 => \N__12850\,
            lcout => \AGNUS_CLK_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;

-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 16 2025 18:12:46

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "U712_TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of U712_TOP
entity U712_TOP is
port (
    CMA : out std_logic_vector(10 downto 0);
    SIZ : in std_logic_vector(1 downto 0);
    DRA : in std_logic_vector(9 downto 0);
    A : in std_logic_vector(20 downto 0);
    RAMENn : out std_logic;
    TSn : in std_logic;
    LMBEn : out std_logic;
    DMA_LATCH_EN : out std_logic;
    CLMBEn : out std_logic;
    AWEn : in std_logic;
    RESETn : in std_logic;
    CLK_EN : out std_logic;
    CASn : out std_logic;
    BANK0 : out std_logic;
    CLK40B_OUT : out std_logic;
    VBENn : out std_logic;
    CUMBEn : out std_logic;
    CLKRAM : out std_logic;
    CLK40D_OUT : out std_logic;
    C3 : in std_logic;
    ASn : out std_logic;
    UUBEn : out std_logic;
    LDSn : out std_logic;
    LATCH_CLK : out std_logic;
    CASUn : in std_logic;
    DRDDIR : out std_logic;
    DBDIR : out std_logic;
    UDSn : out std_logic;
    RnW : in std_logic;
    DRDENn : out std_logic;
    DBENn : out std_logic;
    BANK1 : out std_logic;
    UMBEn : out std_logic;
    RAS0n : in std_logic;
    CUUBEn : out std_logic;
    CRCSn : out std_logic;
    CLLBEn : out std_logic;
    CLK40C_OUT : out std_logic;
    CASLn : in std_logic;
    RAMSPACEn : in std_logic;
    WEn : out std_logic;
    REGENn : out std_logic;
    LLBEn : out std_logic;
    DBRn : in std_logic;
    CLK40_IN : in std_logic;
    REGSPACEn : in std_logic;
    RASn : out std_logic;
    AGNUS_REV : in std_logic;
    TACKn : out std_logic;
    C1 : in std_logic);
end U712_TOP;

-- Architecture of U712_TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of U712_TOP is

signal \N__11850\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11839\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11830\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11821\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11436\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11290\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11272\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11254\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11002\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10983\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10723\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10693\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10691\ : std_logic;
signal \N__10690\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10667\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10661\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10655\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10607\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10574\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10499\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10484\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10469\ : std_logic;
signal \N__10466\ : std_logic;
signal \N__10463\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10457\ : std_logic;
signal \N__10454\ : std_logic;
signal \N__10451\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10408\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10348\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10342\ : std_logic;
signal \N__10339\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10316\ : std_logic;
signal \N__10313\ : std_logic;
signal \N__10310\ : std_logic;
signal \N__10307\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10286\ : std_logic;
signal \N__10283\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10244\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10160\ : std_logic;
signal \N__10157\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10151\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10127\ : std_logic;
signal \N__10124\ : std_logic;
signal \N__10121\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10091\ : std_logic;
signal \N__10088\ : std_logic;
signal \N__10085\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10079\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10019\ : std_logic;
signal \N__10016\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10007\ : std_logic;
signal \N__10004\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9974\ : std_logic;
signal \N__9971\ : std_logic;
signal \N__9970\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9956\ : std_logic;
signal \N__9955\ : std_logic;
signal \N__9952\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9950\ : std_logic;
signal \N__9949\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9797\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9776\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9773\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9770\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9746\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9738\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9735\ : std_logic;
signal \N__9734\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9732\ : std_logic;
signal \N__9731\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9729\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9726\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9723\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9547\ : std_logic;
signal \N__9546\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9437\ : std_logic;
signal \N__9434\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9425\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9407\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9398\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9183\ : std_logic;
signal \N__9180\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9066\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9041\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9014\ : std_logic;
signal \N__9011\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8960\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8936\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8915\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8894\ : std_logic;
signal \N__8885\ : std_logic;
signal \N__8882\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8858\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8801\ : std_logic;
signal \N__8798\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8789\ : std_logic;
signal \N__8786\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8777\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8774\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8725\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8481\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8378\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8342\ : std_logic;
signal \N__8339\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8333\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8331\ : std_logic;
signal \N__8328\ : std_logic;
signal \N__8327\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8256\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8249\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8195\ : std_logic;
signal \N__8192\ : std_logic;
signal \N__8189\ : std_logic;
signal \N__8186\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8180\ : std_logic;
signal \N__8177\ : std_logic;
signal \N__8174\ : std_logic;
signal \N__8171\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8165\ : std_logic;
signal \N__8162\ : std_logic;
signal \N__8159\ : std_logic;
signal \N__8156\ : std_logic;
signal \N__8153\ : std_logic;
signal \N__8150\ : std_logic;
signal \N__8147\ : std_logic;
signal \N__8144\ : std_logic;
signal \N__8141\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8120\ : std_logic;
signal \N__8117\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8111\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8105\ : std_logic;
signal \N__8102\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8096\ : std_logic;
signal \N__8093\ : std_logic;
signal \N__8090\ : std_logic;
signal \N__8087\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8084\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8076\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8051\ : std_logic;
signal \N__8048\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8021\ : std_logic;
signal \N__8018\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7970\ : std_logic;
signal \N__7969\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7957\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7950\ : std_logic;
signal \N__7947\ : std_logic;
signal \N__7944\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7931\ : std_logic;
signal \N__7928\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7923\ : std_logic;
signal \N__7920\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7913\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7875\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7862\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7856\ : std_logic;
signal \N__7851\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7832\ : std_logic;
signal \N__7829\ : std_logic;
signal \N__7826\ : std_logic;
signal \N__7823\ : std_logic;
signal \N__7820\ : std_logic;
signal \N__7817\ : std_logic;
signal \N__7814\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7802\ : std_logic;
signal \N__7799\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7787\ : std_logic;
signal \N__7784\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7772\ : std_logic;
signal \N__7769\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7757\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7721\ : std_logic;
signal \N__7718\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7690\ : std_logic;
signal \N__7687\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7676\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7673\ : std_logic;
signal \N__7658\ : std_logic;
signal \N__7655\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7634\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7622\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7616\ : std_logic;
signal \N__7613\ : std_logic;
signal \N__7610\ : std_logic;
signal \N__7607\ : std_logic;
signal \N__7604\ : std_logic;
signal \N__7601\ : std_logic;
signal \N__7598\ : std_logic;
signal \N__7595\ : std_logic;
signal \N__7592\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7577\ : std_logic;
signal \N__7574\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7565\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7553\ : std_logic;
signal \N__7550\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7520\ : std_logic;
signal \N__7517\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7460\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7430\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7410\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7395\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7349\ : std_logic;
signal \N__7346\ : std_logic;
signal \N__7343\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7337\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7335\ : std_logic;
signal \N__7334\ : std_logic;
signal \N__7331\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7325\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7286\ : std_logic;
signal \N__7283\ : std_logic;
signal \N__7280\ : std_logic;
signal \N__7277\ : std_logic;
signal \N__7274\ : std_logic;
signal \N__7271\ : std_logic;
signal \N__7268\ : std_logic;
signal \N__7265\ : std_logic;
signal \N__7262\ : std_logic;
signal \N__7259\ : std_logic;
signal \N__7256\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7241\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7235\ : std_logic;
signal \N__7232\ : std_logic;
signal \N__7229\ : std_logic;
signal \N__7226\ : std_logic;
signal \N__7223\ : std_logic;
signal \N__7220\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7100\ : std_logic;
signal \N__7097\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7085\ : std_logic;
signal \N__7082\ : std_logic;
signal \N__7079\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7064\ : std_logic;
signal \N__7061\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7026\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6984\ : std_logic;
signal \N__6981\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6956\ : std_logic;
signal \N__6953\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6929\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6917\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6911\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6899\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6893\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6777\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6764\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6708\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6606\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6494\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6446\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6408\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6405\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6393\ : std_logic;
signal \N__6390\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6372\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6336\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6270\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6267\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6213\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6201\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6189\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6154\ : std_logic;
signal \N__6147\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6093\ : std_logic;
signal \N__6090\ : std_logic;
signal \N__6087\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6081\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6057\ : std_logic;
signal \N__6054\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6008\ : std_logic;
signal \N__6005\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5999\ : std_logic;
signal \N__5996\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5904\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5846\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5832\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5778\ : std_logic;
signal \N__5775\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5756\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5744\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5708\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5607\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5600\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5592\ : std_logic;
signal \N__5589\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5333\ : std_logic;
signal \N__5330\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5318\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5235\ : std_logic;
signal \N__5232\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5205\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5184\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5169\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5153\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5129\ : std_logic;
signal \N__5126\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5053\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4986\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4895\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4885\ : std_logic;
signal \N__4882\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4876\ : std_logic;
signal \N__4873\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4831\ : std_logic;
signal \N__4828\ : std_logic;
signal \N__4825\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4770\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4748\ : std_logic;
signal \N__4745\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4724\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4721\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4718\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4688\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4683\ : std_logic;
signal \N__4680\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4637\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4631\ : std_logic;
signal \N__4628\ : std_logic;
signal \N__4625\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4557\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4386\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4378\ : std_logic;
signal \N__4375\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4311\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4288\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4192\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4186\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \CLK40_IN_c\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \CLK80_PLL_i_i\ : std_logic;
signal \U712_CHIP_RAM.N_448_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_459_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_308_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\ : std_logic;
signal \U712_CHIP_RAM.N_416_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_448\ : std_logic;
signal \U712_CHIP_RAM.N_261_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_404_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_413_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_414\ : std_logic;
signal \U712_CHIP_RAM.N_415_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_373_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_373\ : std_logic;
signal \N_48_i\ : std_logic;
signal \RAMSPACEn_c\ : std_logic;
signal \U712_CHIP_RAM.N_355_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\ : std_logic;
signal \TACK_OUTn\ : std_logic;
signal \DBR_SYNCZ0Z_0\ : std_logic;
signal \DBR_SYNCZ0Z_1\ : std_logic;
signal \CLK40_PLL\ : std_logic;
signal \U712_BYTE_ENABLE.N_90\ : std_logic;
signal \CLK40_PLL_g\ : std_logic;
signal \CLK40_PLL_iso_i\ : std_logic;
signal \LATCH_RAM\ : std_logic;
signal \LATCH_CLK_0_i\ : std_logic;
signal \U712_CHIP_RAM.N_296_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_296\ : std_logic;
signal \U712_CHIP_RAM.N_63\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\ : std_logic;
signal \BANK0_c\ : std_logic;
signal \U712_CHIP_RAM.N_404\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\ : std_logic;
signal \A_c_20\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_362\ : std_logic;
signal \U712_CHIP_RAM.N_470\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_344\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0\ : std_logic;
signal \U712_CHIP_RAM.N_344_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_267\ : std_logic;
signal \U712_CHIP_RAM.N_333\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_416\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER_s_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0\ : std_logic;
signal \U712_CHIP_RAM.N_45\ : std_logic;
signal \U712_CHIP_RAM.N_61_cascade_\ : std_logic;
signal \U712_CHIP_RAM.REFRESHZ0\ : std_logic;
signal \U712_CHIP_RAM.N_263\ : std_logic;
signal \U712_CHIP_RAM.N_271\ : std_logic;
signal \U712_CHIP_RAM.N_341_cascade_\ : std_logic;
signal \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_2\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_r_sx_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.CAS_SYNCZ0Z_0\ : std_logic;
signal \U712_CYCLE_TERM.N_286_i_0_0_cascade_\ : std_logic;
signal \U712_CYCLE_TERM.N_286_i_0_en_cascade_\ : std_logic;
signal \RESETn_c_i\ : std_logic;
signal \CPU_TACK\ : std_logic;
signal \U712_CYCLE_TERM.N_286_i_0_en_0\ : std_logic;
signal \DBRn_c\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_0\ : std_logic;
signal \INVU712_REG_SM.DBR_SYNC_1C_net\ : std_logic;
signal \TACK_EN_i_ess\ : std_logic;
signal \N_977_i\ : std_logic;
signal \VBENn_c\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \A_c_6\ : std_logic;
signal \A_c_13\ : std_logic;
signal \A_c_12\ : std_logic;
signal \A_c_5\ : std_logic;
signal \A_c_15\ : std_logic;
signal \A_c_8\ : std_logic;
signal \U712_CHIP_RAM.N_261\ : std_logic;
signal \A_c_11\ : std_logic;
signal \A_c_4\ : std_logic;
signal \U712_CHIP_RAM.N_312\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.N_314\ : std_logic;
signal \U712_CHIP_RAM.N_459\ : std_logic;
signal \U712_CHIP_RAM.N_449\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_\ : std_logic;
signal \RESETn_c\ : std_logic;
signal \U712_CHIP_RAM.N_421\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2\ : std_logic;
signal \U712_CHIP_RAM.N_421_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z20\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_A20C_net\ : std_logic;
signal \U712_CHIP_RAM.N_18\ : std_logic;
signal \U712_CHIP_RAM.N_18_0\ : std_logic;
signal \U712_CHIP_RAM.N_113\ : std_logic;
signal \U712_CHIP_RAM.N_413\ : std_logic;
signal \CLK_EN_c\ : std_logic;
signal \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\ : std_logic;
signal \U712_CHIP_RAM.N_342\ : std_logic;
signal \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\ : std_logic;
signal \AWEn_c\ : std_logic;
signal \DBDIR_c\ : std_logic;
signal \DBRn_c_i\ : std_logic;
signal \DBRn_c_i_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_1\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_4\ : std_logic;
signal \U712_CYCLE_TERM.TACK_STATEZ0Z_0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_5\ : std_logic;
signal \LATCH_REG\ : std_logic;
signal \REG_CPU_CYCLE\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_5C_net\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERc_0_cascade_\ : std_logic;
signal \U712_REG_SM.REG_CPU_CYCLE_e_1\ : std_logic;
signal \A_c_3\ : std_logic;
signal \A_c_10\ : std_logic;
signal \A_c_16\ : std_logic;
signal \A_c_18\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_411_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_\ : std_logic;
signal \U712_CHIP_RAM.N_294\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.N_316_cascade_\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_COUNTER15\ : std_logic;
signal \U712_CHIP_RAM.N_109_i\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERc_0\ : std_logic;
signal \U712_REG_SM.un15_0_i_0_0\ : std_logic;
signal \U712_REG_SM.N_297\ : std_logic;
signal \REG_TACK\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_6\ : std_logic;
signal \REGENn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_4\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_3\ : std_logic;
signal \INVU712_REG_SM.REG_CYCLEC_net\ : std_logic;
signal \U712_REG_SM.DBR_SYNCZ0Z_1\ : std_logic;
signal \INVU712_REG_SM.STATE_COUNTER_2C_net\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\ : std_logic;
signal \A_c_14\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\ : std_logic;
signal \DBENn_c\ : std_logic;
signal \DMA_CYCLE\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lt7\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\ : std_logic;
signal \N_49_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_92\ : std_logic;
signal \N_315\ : std_logic;
signal \U712_REG_SM.N_278_cascade_\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_7\ : std_logic;
signal \U712_REG_SM.N_272\ : std_logic;
signal \U712_REG_SM.N_309\ : std_logic;
signal \U712_REG_SM.N_272_cascade_\ : std_logic;
signal \C3_c\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_0\ : std_logic;
signal \C1_c\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_0\ : std_logic;
signal \U712_REG_SM.LDSn_7_iv_i_0_0\ : std_logic;
signal \U712_REG_SM.N_278\ : std_logic;
signal \ASn_c\ : std_logic;
signal \INVU712_REG_SM.C3_SYNC_0C_net\ : std_logic;
signal \WRITE_CYCLE\ : std_logic;
signal \N_259\ : std_logic;
signal \LDSn_c\ : std_logic;
signal \U712_REG_SM.N_467_cascade_\ : std_logic;
signal \U712_REG_SM.N_371\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\ : std_logic;
signal \CMA_c_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\ : std_logic;
signal \CMA_c_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\ : std_logic;
signal \A_c_7\ : std_logic;
signal \U712_CHIP_RAM.N_329\ : std_logic;
signal \A_c_2\ : std_logic;
signal \A_c_9\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto7_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\ : std_logic;
signal \U712_CHIP_RAM.REFRESH5lto0\ : std_logic;
signal \bfn_12_10_0_\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\ : std_logic;
signal \C1_c_g\ : std_logic;
signal \U712_CHIP_RAM.REFRESH_RST\ : std_logic;
signal \U712_REG_SM.UDSn_7_iv_i_0_0\ : std_logic;
signal \U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1\ : std_logic;
signal \U712_REG_SM.LATCH_REG_0_sqmuxa\ : std_logic;
signal \INVU712_REG_SM.UDSnC_net\ : std_logic;
signal \RAMENn_c\ : std_logic;
signal \TSn_c\ : std_logic;
signal \U712_REG_SM.CYCLE_RUNZ0\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_1\ : std_logic;
signal \RnW_c\ : std_logic;
signal \REG_WRITE_CYCLE\ : std_logic;
signal \INVU712_REG_SM.REG_CYCLE_STARTC_net\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\ : std_logic;
signal \CMA_c_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\ : std_logic;
signal \CMA_c_2\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\ : std_logic;
signal \CMA_c_7\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\ : std_logic;
signal \DRA_c_1\ : std_logic;
signal \DRA_c_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_AZ0Z1\ : std_logic;
signal \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_0\ : std_logic;
signal \U712_REG_SM.N_369\ : std_logic;
signal \UDSn_c\ : std_logic;
signal \U712_REG_SM.STATE_COUNTERZ0Z_2\ : std_logic;
signal \U712_REG_SM.N_465\ : std_logic;
signal \U712_REG_SM.C1_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.REG_CYCLE_STARTZ0\ : std_logic;
signal \U712_REG_SM.C3_SYNCZ0Z_1\ : std_logic;
signal \U712_REG_SM.N_288\ : std_logic;
signal \CASn_c\ : std_logic;
signal \WEn_c\ : std_logic;
signal \RASn_c\ : std_logic;
signal \CRCSn_c\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\ : std_logic;
signal \CMA_c_10\ : std_logic;
signal \A_c_17\ : std_logic;
signal \CMA_c_8\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\ : std_logic;
signal \CMA_c_3\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\ : std_logic;
signal \CMA_c_6\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_sn_N_5_mux\ : std_logic;
signal \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\ : std_logic;
signal \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\ : std_logic;
signal \CMA_c_4\ : std_logic;
signal \A_c_19\ : std_logic;
signal \U712_CHIP_RAM.CMA_5_0_8\ : std_logic;
signal \CMA_c_9\ : std_logic;
signal \CLK80_PLL\ : std_logic;
signal \U712_CHIP_RAM.un1_CMA28_0_i_0\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\ : std_logic;
signal \DRA_c_5\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\ : std_logic;
signal \DRA_c_4\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\ : std_logic;
signal \DRA_c_8\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\ : std_logic;
signal \RAS0n_c\ : std_logic;
signal \DRA_c_9\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\ : std_logic;
signal \DRA_c_6\ : std_logic;
signal \DRA_c_7\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\ : std_logic;
signal \N_50_i\ : std_logic;
signal \CPU_CYCLE\ : std_logic;
signal \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\ : std_logic;
signal \U712_BYTE_ENABLE.N_91_cascade_\ : std_logic;
signal \N_51_i\ : std_logic;
signal \U712_BYTE_ENABLE.N_89\ : std_logic;
signal \N_90_i\ : std_logic;
signal \N_92_i\ : std_logic;
signal \N_91_i\ : std_logic;
signal \SIZ_c_1\ : std_logic;
signal \A_c_1\ : std_logic;
signal \SIZ_c_0\ : std_logic;
signal \A_c_0\ : std_logic;
signal \N_89_i\ : std_logic;
signal \DRA_c_3\ : std_logic;
signal \DRA_c_2\ : std_logic;
signal \AGNUS_REV_c\ : std_logic;
signal \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\ : std_logic;
signal \C3_c_g\ : std_logic;
signal \DBRn_c_i_0_g\ : std_logic;
signal \RESETn_c_i_g\ : std_logic;
signal \REG_CYCLE\ : std_logic;
signal \CASUn_c\ : std_logic;
signal \CASLn_c\ : std_logic;
signal \DRDENn_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DBENn_wire\ : std_logic;
signal \A_wire\ : std_logic_vector(20 downto 0);
signal \CASn_wire\ : std_logic;
signal \DRDDIR_wire\ : std_logic;
signal \C1_wire\ : std_logic;
signal \BANK1_wire\ : std_logic;
signal \DRA_wire\ : std_logic_vector(9 downto 0);
signal \AGNUS_REV_wire\ : std_logic;
signal \RAS0n_wire\ : std_logic;
signal \CMA_wire\ : std_logic_vector(10 downto 0);
signal \UUBEn_wire\ : std_logic;
signal \RAMENn_wire\ : std_logic;
signal \REGSPACEn_wire\ : std_logic;
signal \SIZ_wire\ : std_logic_vector(1 downto 0);
signal \VBENn_wire\ : std_logic;
signal \CASUn_wire\ : std_logic;
signal \DBRn_wire\ : std_logic;
signal \CRCSn_wire\ : std_logic;
signal \LLBEn_wire\ : std_logic;
signal \CASLn_wire\ : std_logic;
signal \TSn_wire\ : std_logic;
signal \RAMSPACEn_wire\ : std_logic;
signal \DMA_LATCH_EN_wire\ : std_logic;
signal \RESETn_wire\ : std_logic;
signal \CLK40_IN_wire\ : std_logic;
signal \RASn_wire\ : std_logic;
signal \BANK0_wire\ : std_logic;
signal \CLK40D_OUT_wire\ : std_logic;
signal \CLKRAM_wire\ : std_logic;
signal \ASn_wire\ : std_logic;
signal \C3_wire\ : std_logic;
signal \CLK40C_OUT_wire\ : std_logic;
signal \DRDENn_wire\ : std_logic;
signal \CLLBEn_wire\ : std_logic;
signal \REGENn_wire\ : std_logic;
signal \CLMBEn_wire\ : std_logic;
signal \WEn_wire\ : std_logic;
signal \DBDIR_wire\ : std_logic;
signal \CUMBEn_wire\ : std_logic;
signal \RnW_wire\ : std_logic;
signal \LMBEn_wire\ : std_logic;
signal \CUUBEn_wire\ : std_logic;
signal \TACKn_wire\ : std_logic;
signal \AWEn_wire\ : std_logic;
signal \UDSn_wire\ : std_logic;
signal \UMBEn_wire\ : std_logic;
signal \CLK_EN_wire\ : std_logic;
signal \LATCH_CLK_wire\ : std_logic;
signal \LDSn_wire\ : std_logic;
signal \CLK40B_OUT_wire\ : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    DBENn <= \DBENn_wire\;
    \A_wire\ <= A;
    CASn <= \CASn_wire\;
    DRDDIR <= \DRDDIR_wire\;
    \C1_wire\ <= C1;
    BANK1 <= \BANK1_wire\;
    \DRA_wire\ <= DRA;
    \AGNUS_REV_wire\ <= AGNUS_REV;
    \RAS0n_wire\ <= RAS0n;
    CMA <= \CMA_wire\;
    UUBEn <= \UUBEn_wire\;
    RAMENn <= \RAMENn_wire\;
    \REGSPACEn_wire\ <= REGSPACEn;
    \SIZ_wire\ <= SIZ;
    VBENn <= \VBENn_wire\;
    \CASUn_wire\ <= CASUn;
    \DBRn_wire\ <= DBRn;
    CRCSn <= \CRCSn_wire\;
    LLBEn <= \LLBEn_wire\;
    \CASLn_wire\ <= CASLn;
    \TSn_wire\ <= TSn;
    \RAMSPACEn_wire\ <= RAMSPACEn;
    DMA_LATCH_EN <= \DMA_LATCH_EN_wire\;
    \RESETn_wire\ <= RESETn;
    \CLK40_IN_wire\ <= CLK40_IN;
    RASn <= \RASn_wire\;
    BANK0 <= \BANK0_wire\;
    CLK40D_OUT <= \CLK40D_OUT_wire\;
    CLKRAM <= \CLKRAM_wire\;
    ASn <= \ASn_wire\;
    \C3_wire\ <= C3;
    CLK40C_OUT <= \CLK40C_OUT_wire\;
    DRDENn <= \DRDENn_wire\;
    CLLBEn <= \CLLBEn_wire\;
    REGENn <= \REGENn_wire\;
    CLMBEn <= \CLMBEn_wire\;
    WEn <= \WEn_wire\;
    DBDIR <= \DBDIR_wire\;
    CUMBEn <= \CUMBEn_wire\;
    \RnW_wire\ <= RnW;
    LMBEn <= \LMBEn_wire\;
    CUUBEn <= \CUUBEn_wire\;
    TACKn <= \TACKn_wire\;
    \AWEn_wire\ <= AWEn;
    UDSn <= \UDSn_wire\;
    UMBEn <= \UMBEn_wire\;
    CLK_EN <= \CLK_EN_wire\;
    LATCH_CLK <= \LATCH_CLK_wire\;
    LDSn <= \LDSn_wire\;
    CLK40B_OUT <= \CLK40B_OUT_wire\;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "DELAY",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "011",
            DIVF => "0000001",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => \CLK40_PLL\,
            REFERENCECLK => \N__4061\,
            RESETB => \N__4901\,
            BYPASS => '0',
            PLLOUTCOREA => OPEN,
            SDI => '0',
            PLLOUTGLOBALB => OPEN,
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => '0',
            PLLOUTGLOBALA => \CLK80_PLL\,
            SCLK => '0'
        );

    \DBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11850\,
            DIN => \N__11849\,
            DOUT => \N__11848\,
            PACKAGEPIN => \DBENn_wire\
        );

    \DBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11850\,
            PADOUT => \N__11849\,
            PADIN => \N__11848\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7052\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11841\,
            DIN => \N__11840\,
            DOUT => \N__11839\,
            PACKAGEPIN => \A_wire\(2)
        );

    \A_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11841\,
            PADOUT => \N__11840\,
            PADIN => \N__11839\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11832\,
            DIN => \N__11831\,
            DOUT => \N__11830\,
            PACKAGEPIN => \CASn_wire\
        );

    \CASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11832\,
            PADOUT => \N__11831\,
            PADIN => \N__11830\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8198\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11823\,
            DIN => \N__11822\,
            DOUT => \N__11821\,
            PACKAGEPIN => \DRDDIR_wire\
        );

    \DRDDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11823\,
            PADOUT => \N__11822\,
            PADIN => \N__11821\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7241\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11814\,
            DIN => \N__11813\,
            DOUT => \N__11812\,
            PACKAGEPIN => \C1_wire\
        );

    \C1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11814\,
            PADOUT => \N__11813\,
            PADIN => \N__11812\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11805\,
            DIN => \N__11804\,
            DOUT => \N__11803\,
            PACKAGEPIN => \BANK1_wire\
        );

    \BANK1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11805\,
            PADOUT => \N__11804\,
            PADIN => \N__11803\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11796\,
            DIN => \N__11795\,
            DOUT => \N__11794\,
            PACKAGEPIN => \DRA_wire\(3)
        );

    \DRA_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11796\,
            PADOUT => \N__11795\,
            PADIN => \N__11794\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AGNUS_REV_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11787\,
            DIN => \N__11786\,
            DOUT => \N__11785\,
            PACKAGEPIN => \AGNUS_REV_wire\
        );

    \AGNUS_REV_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11787\,
            PADOUT => \N__11786\,
            PADIN => \N__11785\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AGNUS_REV_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAS0n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11778\,
            DIN => \N__11777\,
            DOUT => \N__11776\,
            PACKAGEPIN => \RAS0n_wire\
        );

    \RAS0n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11778\,
            PADOUT => \N__11777\,
            PADIN => \N__11776\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAS0n_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11769\,
            DIN => \N__11768\,
            DOUT => \N__11767\,
            PACKAGEPIN => \A_wire\(7)
        );

    \A_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11769\,
            PADOUT => \N__11768\,
            PADIN => \N__11767\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11760\,
            DIN => \N__11759\,
            DOUT => \N__11758\,
            PACKAGEPIN => \CMA_wire\(7)
        );

    \CMA_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11760\,
            PADOUT => \N__11759\,
            PADIN => \N__11758\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11751\,
            DIN => \N__11750\,
            DOUT => \N__11749\,
            PACKAGEPIN => \UUBEn_wire\
        );

    \UUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11751\,
            PADOUT => \N__11750\,
            PADIN => \N__11749\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10436\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11742\,
            DIN => \N__11741\,
            DOUT => \N__11740\,
            PACKAGEPIN => \DRA_wire\(9)
        );

    \DRA_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11742\,
            PADOUT => \N__11741\,
            PADIN => \N__11740\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11733\,
            DIN => \N__11732\,
            DOUT => \N__11731\,
            PACKAGEPIN => \RAMENn_wire\
        );

    \RAMENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11733\,
            PADOUT => \N__11732\,
            PADIN => \N__11731\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8051\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11724\,
            DIN => \N__11723\,
            DOUT => \N__11722\,
            PACKAGEPIN => \REGSPACEn_wire\
        );

    \REGSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11724\,
            PADOUT => \N__11723\,
            PADIN => \N__11722\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMENn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11715\,
            DIN => \N__11714\,
            DOUT => \N__11713\,
            PACKAGEPIN => \SIZ_wire\(0)
        );

    \SIZ_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11715\,
            PADOUT => \N__11714\,
            PADIN => \N__11713\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \VBENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11706\,
            DIN => \N__11705\,
            DOUT => \N__11704\,
            PACKAGEPIN => \VBENn_wire\
        );

    \VBENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11706\,
            PADOUT => \N__11705\,
            PADIN => \N__11704\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4919\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASUn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11697\,
            DIN => \N__11696\,
            DOUT => \N__11695\,
            PACKAGEPIN => \CASUn_wire\
        );

    \CASUn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11697\,
            PADOUT => \N__11696\,
            PADIN => \N__11695\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASUn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11688\,
            DIN => \N__11687\,
            DOUT => \N__11686\,
            PACKAGEPIN => \A_wire\(4)
        );

    \A_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11688\,
            PADOUT => \N__11687\,
            PADIN => \N__11686\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11679\,
            DIN => \N__11678\,
            DOUT => \N__11677\,
            PACKAGEPIN => \CMA_wire\(0)
        );

    \CMA_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11679\,
            PADOUT => \N__11678\,
            PADIN => \N__11677\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7841\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBRn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11670\,
            DIN => \N__11669\,
            DOUT => \N__11668\,
            PACKAGEPIN => \DBRn_wire\
        );

    \DBRn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11670\,
            PADOUT => \N__11669\,
            PADIN => \N__11668\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DBRn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CRCSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11661\,
            DIN => \N__11660\,
            DOUT => \N__11659\,
            PACKAGEPIN => \CRCSn_wire\
        );

    \CRCSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11661\,
            PADOUT => \N__11660\,
            PADIN => \N__11659\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9209\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11652\,
            DIN => \N__11651\,
            DOUT => \N__11650\,
            PACKAGEPIN => \A_wire\(12)
        );

    \A_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11652\,
            PADOUT => \N__11651\,
            PADIN => \N__11650\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_12\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11643\,
            DIN => \N__11642\,
            DOUT => \N__11641\,
            PACKAGEPIN => \LLBEn_wire\
        );

    \LLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11643\,
            PADOUT => \N__11642\,
            PADIN => \N__11641\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10469\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CASLn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11634\,
            DIN => \N__11633\,
            DOUT => \N__11632\,
            PACKAGEPIN => \CASLn_wire\
        );

    \CASLn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11634\,
            PADOUT => \N__11633\,
            PADIN => \N__11632\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CASLn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TSn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11625\,
            DIN => \N__11624\,
            DOUT => \N__11623\,
            PACKAGEPIN => \TSn_wire\
        );

    \TSn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11625\,
            PADOUT => \N__11624\,
            PADIN => \N__11623\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TSn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RAMSPACEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11616\,
            DIN => \N__11615\,
            DOUT => \N__11614\,
            PACKAGEPIN => \RAMSPACEn_wire\
        );

    \RAMSPACEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11616\,
            PADOUT => \N__11615\,
            PADIN => \N__11614\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RAMSPACEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11607\,
            DIN => \N__11606\,
            DOUT => \N__11605\,
            PACKAGEPIN => \A_wire\(18)
        );

    \A_ibuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11607\,
            PADOUT => \N__11606\,
            PADIN => \N__11605\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_18\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11598\,
            DIN => \N__11597\,
            DOUT => \N__11596\,
            PACKAGEPIN => \A_wire\(9)
        );

    \A_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11598\,
            PADOUT => \N__11597\,
            PADIN => \N__11596\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DMA_LATCH_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11589\,
            DIN => \N__11588\,
            DOUT => \N__11587\,
            PACKAGEPIN => \DMA_LATCH_EN_wire\
        );

    \DMA_LATCH_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11589\,
            PADOUT => \N__11588\,
            PADIN => \N__11587\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11580\,
            DIN => \N__11579\,
            DOUT => \N__11578\,
            PACKAGEPIN => \DRA_wire\(7)
        );

    \DRA_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11580\,
            PADOUT => \N__11579\,
            PADIN => \N__11578\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11571\,
            DIN => \N__11570\,
            DOUT => \N__11569\,
            PACKAGEPIN => \A_wire\(15)
        );

    \A_ibuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11571\,
            PADOUT => \N__11570\,
            PADIN => \N__11569\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_15\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RESETn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11562\,
            DIN => \N__11561\,
            DOUT => \N__11560\,
            PACKAGEPIN => \RESETn_wire\
        );

    \RESETn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11562\,
            PADOUT => \N__11561\,
            PADIN => \N__11560\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RESETn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11553\,
            DIN => \N__11552\,
            DOUT => \N__11551\,
            PACKAGEPIN => \A_wire\(3)
        );

    \A_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11553\,
            PADOUT => \N__11552\,
            PADIN => \N__11551\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40_IN_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11544\,
            DIN => \N__11543\,
            DOUT => \N__11542\,
            PACKAGEPIN => \CLK40_IN_wire\
        );

    \CLK40_IN_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11544\,
            PADOUT => \N__11543\,
            PADIN => \N__11542\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \CLK40_IN_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11535\,
            DIN => \N__11534\,
            DOUT => \N__11533\,
            PACKAGEPIN => \RASn_wire\
        );

    \RASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11535\,
            PADOUT => \N__11534\,
            PADIN => \N__11533\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9227\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \BANK0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11526\,
            DIN => \N__11525\,
            DOUT => \N__11524\,
            PACKAGEPIN => \BANK0_wire\
        );

    \BANK0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11526\,
            PADOUT => \N__11525\,
            PADIN => \N__11524\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4475\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40D_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11517\,
            DIN => \N__11516\,
            DOUT => \N__11515\,
            PACKAGEPIN => \CLK40D_OUT_wire\
        );

    \CLK40D_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11517\,
            PADOUT => \N__11516\,
            PADIN => \N__11515\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4216\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLKRAM_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11508\,
            DIN => \N__11507\,
            DOUT => \N__11506\,
            PACKAGEPIN => \CLKRAM_wire\
        );

    \CLKRAM_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11508\,
            PADOUT => \N__11507\,
            PADIN => \N__11506\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4091\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11499\,
            DIN => \N__11498\,
            DOUT => \N__11497\,
            PACKAGEPIN => \DRA_wire\(0)
        );

    \DRA_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11499\,
            PADOUT => \N__11498\,
            PADIN => \N__11497\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ASn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11490\,
            DIN => \N__11489\,
            DOUT => \N__11488\,
            PACKAGEPIN => \ASn_wire\
        );

    \ASn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11490\,
            PADOUT => \N__11489\,
            PADIN => \N__11488\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7457\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11481\,
            DIN => \N__11480\,
            DOUT => \N__11479\,
            PACKAGEPIN => \CMA_wire\(3)
        );

    \CMA_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11481\,
            PADOUT => \N__11480\,
            PADIN => \N__11479\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8822\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11472\,
            DIN => \N__11471\,
            DOUT => \N__11470\,
            PACKAGEPIN => \A_wire\(20)
        );

    \A_ibuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11472\,
            PADOUT => \N__11471\,
            PADIN => \N__11470\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_20\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \C3_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11463\,
            DIN => \N__11462\,
            DOUT => \N__11461\,
            PACKAGEPIN => \C3_wire\
        );

    \C3_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11463\,
            PADOUT => \N__11462\,
            PADIN => \N__11461\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \C3_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11454\,
            DIN => \N__11453\,
            DOUT => \N__11452\,
            PACKAGEPIN => \DRA_wire\(5)
        );

    \DRA_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11454\,
            PADOUT => \N__11453\,
            PADIN => \N__11452\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11445\,
            DIN => \N__11444\,
            DOUT => \N__11443\,
            PACKAGEPIN => \A_wire\(0)
        );

    \A_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11445\,
            PADOUT => \N__11444\,
            PADIN => \N__11443\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_0\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11436\,
            DIN => \N__11435\,
            DOUT => \N__11434\,
            PACKAGEPIN => \CMA_wire\(10)
        );

    \CMA_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11436\,
            PADOUT => \N__11435\,
            PADIN => \N__11434\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8885\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11427\,
            DIN => \N__11426\,
            DOUT => \N__11425\,
            PACKAGEPIN => \A_wire\(13)
        );

    \A_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11427\,
            PADOUT => \N__11426\,
            PADIN => \N__11425\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_13\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40C_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11418\,
            DIN => \N__11417\,
            DOUT => \N__11416\,
            PACKAGEPIN => \CLK40C_OUT_wire\
        );

    \CLK40C_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11418\,
            PADOUT => \N__11417\,
            PADIN => \N__11416\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4204\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11409\,
            DIN => \N__11408\,
            DOUT => \N__11407\,
            PACKAGEPIN => \CMA_wire\(4)
        );

    \CMA_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11409\,
            PADOUT => \N__11408\,
            PADIN => \N__11407\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8687\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRDENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11400\,
            DIN => \N__11399\,
            DOUT => \N__11398\,
            PACKAGEPIN => \DRDENn_wire\
        );

    \DRDENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11400\,
            PADOUT => \N__11399\,
            PADIN => \N__11398\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10715\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLLBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11391\,
            DIN => \N__11390\,
            DOUT => \N__11389\,
            PACKAGEPIN => \CLLBEn_wire\
        );

    \CLLBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11391\,
            PADOUT => \N__11390\,
            PADIN => \N__11389\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4142\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11382\,
            DIN => \N__11381\,
            DOUT => \N__11380\,
            PACKAGEPIN => \CMA_wire\(9)
        );

    \CMA_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11382\,
            PADOUT => \N__11381\,
            PADIN => \N__11380\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8615\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \REGENn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11373\,
            DIN => \N__11372\,
            DOUT => \N__11371\,
            PACKAGEPIN => \REGENn_wire\
        );

    \REGENn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11373\,
            PADOUT => \N__11372\,
            PADIN => \N__11371\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6818\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11364\,
            DIN => \N__11363\,
            DOUT => \N__11362\,
            PACKAGEPIN => \A_wire\(19)
        );

    \A_ibuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11364\,
            PADOUT => \N__11363\,
            PADIN => \N__11362\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_19\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11355\,
            DIN => \N__11354\,
            DOUT => \N__11353\,
            PACKAGEPIN => \A_wire\(8)
        );

    \A_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11355\,
            PADOUT => \N__11354\,
            PADIN => \N__11353\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11346\,
            DIN => \N__11345\,
            DOUT => \N__11344\,
            PACKAGEPIN => \CLMBEn_wire\
        );

    \CLMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11346\,
            PADOUT => \N__11345\,
            PADIN => \N__11344\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6929\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \WEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11337\,
            DIN => \N__11336\,
            DOUT => \N__11335\,
            PACKAGEPIN => \WEn_wire\
        );

    \WEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11337\,
            PADOUT => \N__11336\,
            PADIN => \N__11335\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DBDIR_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11328\,
            DIN => \N__11327\,
            DOUT => \N__11326\,
            PACKAGEPIN => \DBDIR_wire\
        );

    \DBDIR_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11328\,
            PADOUT => \N__11327\,
            PADIN => \N__11326\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5492\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11319\,
            DIN => \N__11318\,
            DOUT => \N__11317\,
            PACKAGEPIN => \CUMBEn_wire\
        );

    \CUMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11319\,
            PADOUT => \N__11318\,
            PADIN => \N__11317\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11310\,
            DIN => \N__11309\,
            DOUT => \N__11308\,
            PACKAGEPIN => \DRA_wire\(6)
        );

    \DRA_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11310\,
            PADOUT => \N__11309\,
            PADIN => \N__11308\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11301\,
            DIN => \N__11300\,
            DOUT => \N__11299\,
            PACKAGEPIN => \A_wire\(5)
        );

    \A_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11301\,
            PADOUT => \N__11300\,
            PADIN => \N__11299\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \RnW_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11292\,
            DIN => \N__11291\,
            DOUT => \N__11290\,
            PACKAGEPIN => \RnW_wire\
        );

    \RnW_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11292\,
            PADOUT => \N__11291\,
            PADIN => \N__11290\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \RnW_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11283\,
            DIN => \N__11282\,
            DOUT => \N__11281\,
            PACKAGEPIN => \A_wire\(16)
        );

    \A_ibuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11283\,
            PADOUT => \N__11282\,
            PADIN => \N__11281\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_16\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11274\,
            DIN => \N__11273\,
            DOUT => \N__11272\,
            PACKAGEPIN => \CMA_wire\(1)
        );

    \CMA_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11274\,
            PADOUT => \N__11273\,
            PADIN => \N__11272\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7298\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11265\,
            DIN => \N__11264\,
            DOUT => \N__11263\,
            PACKAGEPIN => \LMBEn_wire\
        );

    \LMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11265\,
            PADOUT => \N__11264\,
            PADIN => \N__11263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10454\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11256\,
            DIN => \N__11255\,
            DOUT => \N__11254\,
            PACKAGEPIN => \A_wire\(11)
        );

    \A_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11256\,
            PADOUT => \N__11255\,
            PADIN => \N__11254\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_11\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CUUBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11247\,
            DIN => \N__11246\,
            DOUT => \N__11245\,
            PACKAGEPIN => \CUUBEn_wire\
        );

    \CUUBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11247\,
            PADOUT => \N__11246\,
            PADIN => \N__11245\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10496\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TACKn_obuft_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11238\,
            DIN => \N__11237\,
            DOUT => \N__11236\,
            PACKAGEPIN => \TACKn_wire\
        );

    \TACKn_obuft_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "101001"
        )
    port map (
            PADOEN => \N__11238\,
            PADOUT => \N__11237\,
            PADIN => \N__11236\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__4940\,
            DIN0 => OPEN,
            DOUT0 => \N__4364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11229\,
            DIN => \N__11228\,
            DOUT => \N__11227\,
            PACKAGEPIN => \CMA_wire\(2)
        );

    \CMA_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11229\,
            PADOUT => \N__11228\,
            PADIN => \N__11227\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7817\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11220\,
            DIN => \N__11219\,
            DOUT => \N__11218\,
            PACKAGEPIN => \DRA_wire\(4)
        );

    \DRA_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11220\,
            PADOUT => \N__11219\,
            PADIN => \N__11218\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11211\,
            DIN => \N__11210\,
            DOUT => \N__11209\,
            PACKAGEPIN => \A_wire\(14)
        );

    \A_ibuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11211\,
            PADOUT => \N__11210\,
            PADIN => \N__11209\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_14\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11202\,
            DIN => \N__11201\,
            DOUT => \N__11200\,
            PACKAGEPIN => \CMA_wire\(8)
        );

    \CMA_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11202\,
            PADOUT => \N__11201\,
            PADIN => \N__11200\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8852\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \AWEn_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11193\,
            DIN => \N__11192\,
            DOUT => \N__11191\,
            PACKAGEPIN => \AWEn_wire\
        );

    \AWEn_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11193\,
            PADOUT => \N__11192\,
            PADIN => \N__11191\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \AWEn_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11184\,
            DIN => \N__11183\,
            DOUT => \N__11182\,
            PACKAGEPIN => \DRA_wire\(1)
        );

    \DRA_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11184\,
            PADOUT => \N__11183\,
            PADIN => \N__11182\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11175\,
            DIN => \N__11174\,
            DOUT => \N__11173\,
            PACKAGEPIN => \A_wire\(17)
        );

    \A_ibuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11175\,
            PADOUT => \N__11174\,
            PADIN => \N__11173\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_17\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11166\,
            DIN => \N__11165\,
            DOUT => \N__11164\,
            PACKAGEPIN => \A_wire\(1)
        );

    \A_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11166\,
            PADOUT => \N__11165\,
            PADIN => \N__11164\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11157\,
            DIN => \N__11156\,
            DOUT => \N__11155\,
            PACKAGEPIN => \CMA_wire\(5)
        );

    \CMA_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11157\,
            PADOUT => \N__11156\,
            PADIN => \N__11155\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7277\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11148\,
            DIN => \N__11147\,
            DOUT => \N__11146\,
            PACKAGEPIN => \UDSn_wire\
        );

    \UDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11148\,
            PADOUT => \N__11147\,
            PADIN => \N__11146\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8441\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \UMBEn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11139\,
            DIN => \N__11138\,
            DOUT => \N__11137\,
            PACKAGEPIN => \UMBEn_wire\
        );

    \UMBEn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11139\,
            PADOUT => \N__11138\,
            PADIN => \N__11137\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10094\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK_EN_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11130\,
            DIN => \N__11129\,
            DOUT => \N__11128\,
            PACKAGEPIN => \CLK_EN_wire\
        );

    \CLK_EN_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11130\,
            PADOUT => \N__11129\,
            PADIN => \N__11128\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5582\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11121\,
            DIN => \N__11120\,
            DOUT => \N__11119\,
            PACKAGEPIN => \DRA_wire\(2)
        );

    \DRA_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11121\,
            PADOUT => \N__11120\,
            PADIN => \N__11119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11112\,
            DIN => \N__11111\,
            DOUT => \N__11110\,
            PACKAGEPIN => \A_wire\(6)
        );

    \A_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11112\,
            PADOUT => \N__11111\,
            PADIN => \N__11110\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CMA_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11103\,
            DIN => \N__11102\,
            DOUT => \N__11101\,
            PACKAGEPIN => \CMA_wire\(6)
        );

    \CMA_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11103\,
            PADOUT => \N__11102\,
            PADIN => \N__11101\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8801\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DRA_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11094\,
            DIN => \N__11093\,
            DOUT => \N__11092\,
            PACKAGEPIN => \DRA_wire\(8)
        );

    \DRA_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11094\,
            PADOUT => \N__11093\,
            PADIN => \N__11092\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DRA_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \A_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11085\,
            DIN => \N__11084\,
            DOUT => \N__11083\,
            PACKAGEPIN => \A_wire\(10)
        );

    \A_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11085\,
            PADOUT => \N__11084\,
            PADIN => \N__11083\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \A_c_10\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LATCH_CLK_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11076\,
            DIN => \N__11075\,
            DOUT => \N__11074\,
            PACKAGEPIN => \LATCH_CLK_wire\
        );

    \LATCH_CLK_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11076\,
            PADOUT => \N__11075\,
            PADIN => \N__11074\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4424\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LDSn_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11067\,
            DIN => \N__11066\,
            DOUT => \N__11065\,
            PACKAGEPIN => \LDSn_wire\
        );

    \LDSn_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11067\,
            PADOUT => \N__11066\,
            PADIN => \N__11065\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \CLK40B_OUT_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11058\,
            DIN => \N__11057\,
            DOUT => \N__11056\,
            PACKAGEPIN => \CLK40B_OUT_wire\
        );

    \CLK40B_OUT_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__11058\,
            PADOUT => \N__11057\,
            PADIN => \N__11056\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4217\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \SIZ_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__11049\,
            DIN => \N__11048\,
            DOUT => \N__11047\,
            PACKAGEPIN => \SIZ_wire\(1)
        );

    \SIZ_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__11049\,
            PADOUT => \N__11048\,
            PADIN => \N__11047\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \SIZ_c_1\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2684\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11024\
        );

    \I__2683\ : InMux
    port map (
            O => \N__11029\,
            I => \N__11021\
        );

    \I__2682\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11018\
        );

    \I__2681\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11015\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__11024\,
            I => \N__11009\
        );

    \I__2679\ : LocalMux
    port map (
            O => \N__11021\,
            I => \N__11004\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11018\,
            I => \N__10996\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__11015\,
            I => \N__10984\
        );

    \I__2676\ : SRMux
    port map (
            O => \N__11014\,
            I => \N__10901\
        );

    \I__2675\ : SRMux
    port map (
            O => \N__11013\,
            I => \N__10901\
        );

    \I__2674\ : SRMux
    port map (
            O => \N__11012\,
            I => \N__10901\
        );

    \I__2673\ : Glb2LocalMux
    port map (
            O => \N__11009\,
            I => \N__10901\
        );

    \I__2672\ : SRMux
    port map (
            O => \N__11008\,
            I => \N__10901\
        );

    \I__2671\ : SRMux
    port map (
            O => \N__11007\,
            I => \N__10901\
        );

    \I__2670\ : Glb2LocalMux
    port map (
            O => \N__11004\,
            I => \N__10901\
        );

    \I__2669\ : SRMux
    port map (
            O => \N__11003\,
            I => \N__10901\
        );

    \I__2668\ : SRMux
    port map (
            O => \N__11002\,
            I => \N__10901\
        );

    \I__2667\ : SRMux
    port map (
            O => \N__11001\,
            I => \N__10901\
        );

    \I__2666\ : SRMux
    port map (
            O => \N__11000\,
            I => \N__10901\
        );

    \I__2665\ : SRMux
    port map (
            O => \N__10999\,
            I => \N__10901\
        );

    \I__2664\ : Glb2LocalMux
    port map (
            O => \N__10996\,
            I => \N__10901\
        );

    \I__2663\ : SRMux
    port map (
            O => \N__10995\,
            I => \N__10901\
        );

    \I__2662\ : SRMux
    port map (
            O => \N__10994\,
            I => \N__10901\
        );

    \I__2661\ : SRMux
    port map (
            O => \N__10993\,
            I => \N__10901\
        );

    \I__2660\ : SRMux
    port map (
            O => \N__10992\,
            I => \N__10901\
        );

    \I__2659\ : SRMux
    port map (
            O => \N__10991\,
            I => \N__10901\
        );

    \I__2658\ : SRMux
    port map (
            O => \N__10990\,
            I => \N__10901\
        );

    \I__2657\ : SRMux
    port map (
            O => \N__10989\,
            I => \N__10901\
        );

    \I__2656\ : SRMux
    port map (
            O => \N__10988\,
            I => \N__10901\
        );

    \I__2655\ : SRMux
    port map (
            O => \N__10987\,
            I => \N__10901\
        );

    \I__2654\ : Glb2LocalMux
    port map (
            O => \N__10984\,
            I => \N__10901\
        );

    \I__2653\ : SRMux
    port map (
            O => \N__10983\,
            I => \N__10901\
        );

    \I__2652\ : SRMux
    port map (
            O => \N__10982\,
            I => \N__10901\
        );

    \I__2651\ : SRMux
    port map (
            O => \N__10981\,
            I => \N__10901\
        );

    \I__2650\ : SRMux
    port map (
            O => \N__10980\,
            I => \N__10901\
        );

    \I__2649\ : SRMux
    port map (
            O => \N__10979\,
            I => \N__10901\
        );

    \I__2648\ : SRMux
    port map (
            O => \N__10978\,
            I => \N__10901\
        );

    \I__2647\ : SRMux
    port map (
            O => \N__10977\,
            I => \N__10901\
        );

    \I__2646\ : SRMux
    port map (
            O => \N__10976\,
            I => \N__10901\
        );

    \I__2645\ : SRMux
    port map (
            O => \N__10975\,
            I => \N__10901\
        );

    \I__2644\ : SRMux
    port map (
            O => \N__10974\,
            I => \N__10901\
        );

    \I__2643\ : SRMux
    port map (
            O => \N__10973\,
            I => \N__10901\
        );

    \I__2642\ : SRMux
    port map (
            O => \N__10972\,
            I => \N__10901\
        );

    \I__2641\ : GlobalMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__2640\ : gio2CtrlBuf
    port map (
            O => \N__10898\,
            I => \RESETn_c_i_g\
        );

    \I__2639\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__10889\,
            I => \N__10886\
        );

    \I__2636\ : Span4Mux_h
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__2635\ : Span4Mux_h
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10876\
        );

    \I__2633\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10873\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__10876\,
            I => \REG_CYCLE\
        );

    \I__2631\ : LocalMux
    port map (
            O => \N__10873\,
            I => \REG_CYCLE\
        );

    \I__2630\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10865\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10861\
        );

    \I__2628\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10858\
        );

    \I__2627\ : Span4Mux_v
    port map (
            O => \N__10861\,
            I => \N__10854\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__10858\,
            I => \N__10851\
        );

    \I__2625\ : InMux
    port map (
            O => \N__10857\,
            I => \N__10848\
        );

    \I__2624\ : Span4Mux_h
    port map (
            O => \N__10854\,
            I => \N__10841\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__10851\,
            I => \N__10841\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__10848\,
            I => \N__10841\
        );

    \I__2621\ : Span4Mux_v
    port map (
            O => \N__10841\,
            I => \N__10838\
        );

    \I__2620\ : Span4Mux_h
    port map (
            O => \N__10838\,
            I => \N__10833\
        );

    \I__2619\ : InMux
    port map (
            O => \N__10837\,
            I => \N__10829\
        );

    \I__2618\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10826\
        );

    \I__2617\ : Span4Mux_h
    port map (
            O => \N__10833\,
            I => \N__10823\
        );

    \I__2616\ : InMux
    port map (
            O => \N__10832\,
            I => \N__10820\
        );

    \I__2615\ : LocalMux
    port map (
            O => \N__10829\,
            I => \N__10817\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__10826\,
            I => \N__10814\
        );

    \I__2613\ : Span4Mux_h
    port map (
            O => \N__10823\,
            I => \N__10809\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10809\
        );

    \I__2611\ : Span12Mux_h
    port map (
            O => \N__10817\,
            I => \N__10806\
        );

    \I__2610\ : Span12Mux_v
    port map (
            O => \N__10814\,
            I => \N__10803\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__10809\,
            I => \N__10800\
        );

    \I__2608\ : Span12Mux_v
    port map (
            O => \N__10806\,
            I => \N__10797\
        );

    \I__2607\ : Span12Mux_h
    port map (
            O => \N__10803\,
            I => \N__10794\
        );

    \I__2606\ : Span4Mux_v
    port map (
            O => \N__10800\,
            I => \N__10791\
        );

    \I__2605\ : Odrv12
    port map (
            O => \N__10797\,
            I => \CASUn_c\
        );

    \I__2604\ : Odrv12
    port map (
            O => \N__10794\,
            I => \CASUn_c\
        );

    \I__2603\ : Odrv4
    port map (
            O => \N__10791\,
            I => \CASUn_c\
        );

    \I__2602\ : InMux
    port map (
            O => \N__10784\,
            I => \N__10779\
        );

    \I__2601\ : InMux
    port map (
            O => \N__10783\,
            I => \N__10776\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__10782\,
            I => \N__10772\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__10779\,
            I => \N__10767\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__10776\,
            I => \N__10767\
        );

    \I__2597\ : InMux
    port map (
            O => \N__10775\,
            I => \N__10764\
        );

    \I__2596\ : InMux
    port map (
            O => \N__10772\,
            I => \N__10760\
        );

    \I__2595\ : Span4Mux_v
    port map (
            O => \N__10767\,
            I => \N__10755\
        );

    \I__2594\ : LocalMux
    port map (
            O => \N__10764\,
            I => \N__10755\
        );

    \I__2593\ : InMux
    port map (
            O => \N__10763\,
            I => \N__10752\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__10760\,
            I => \N__10749\
        );

    \I__2591\ : Span4Mux_h
    port map (
            O => \N__10755\,
            I => \N__10744\
        );

    \I__2590\ : LocalMux
    port map (
            O => \N__10752\,
            I => \N__10744\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__10749\,
            I => \N__10741\
        );

    \I__2588\ : Sp12to4
    port map (
            O => \N__10744\,
            I => \N__10737\
        );

    \I__2587\ : Sp12to4
    port map (
            O => \N__10741\,
            I => \N__10734\
        );

    \I__2586\ : InMux
    port map (
            O => \N__10740\,
            I => \N__10731\
        );

    \I__2585\ : Span12Mux_v
    port map (
            O => \N__10737\,
            I => \N__10728\
        );

    \I__2584\ : Span12Mux_h
    port map (
            O => \N__10734\,
            I => \N__10723\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__10731\,
            I => \N__10723\
        );

    \I__2582\ : Span12Mux_h
    port map (
            O => \N__10728\,
            I => \N__10718\
        );

    \I__2581\ : Span12Mux_v
    port map (
            O => \N__10723\,
            I => \N__10718\
        );

    \I__2580\ : Odrv12
    port map (
            O => \N__10718\,
            I => \CASLn_c\
        );

    \I__2579\ : IoInMux
    port map (
            O => \N__10715\,
            I => \N__10712\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__10712\,
            I => \N__10709\
        );

    \I__2577\ : Span4Mux_s3_v
    port map (
            O => \N__10709\,
            I => \N__10706\
        );

    \I__2576\ : Span4Mux_v
    port map (
            O => \N__10706\,
            I => \N__10703\
        );

    \I__2575\ : Sp12to4
    port map (
            O => \N__10703\,
            I => \N__10700\
        );

    \I__2574\ : Odrv12
    port map (
            O => \N__10700\,
            I => \DRDENn_c\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__10697\,
            I => \N__10694\
        );

    \I__2572\ : InMux
    port map (
            O => \N__10694\,
            I => \N__10687\
        );

    \I__2571\ : CascadeMux
    port map (
            O => \N__10693\,
            I => \N__10683\
        );

    \I__2570\ : CascadeMux
    port map (
            O => \N__10692\,
            I => \N__10680\
        );

    \I__2569\ : CascadeMux
    port map (
            O => \N__10691\,
            I => \N__10675\
        );

    \I__2568\ : InMux
    port map (
            O => \N__10690\,
            I => \N__10667\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__10687\,
            I => \N__10664\
        );

    \I__2566\ : InMux
    port map (
            O => \N__10686\,
            I => \N__10661\
        );

    \I__2565\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10656\
        );

    \I__2564\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10656\
        );

    \I__2563\ : InMux
    port map (
            O => \N__10679\,
            I => \N__10651\
        );

    \I__2562\ : InMux
    port map (
            O => \N__10678\,
            I => \N__10648\
        );

    \I__2561\ : InMux
    port map (
            O => \N__10675\,
            I => \N__10642\
        );

    \I__2560\ : CascadeMux
    port map (
            O => \N__10674\,
            I => \N__10636\
        );

    \I__2559\ : InMux
    port map (
            O => \N__10673\,
            I => \N__10626\
        );

    \I__2558\ : InMux
    port map (
            O => \N__10672\,
            I => \N__10626\
        );

    \I__2557\ : InMux
    port map (
            O => \N__10671\,
            I => \N__10626\
        );

    \I__2556\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10626\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__10667\,
            I => \N__10617\
        );

    \I__2554\ : Span4Mux_h
    port map (
            O => \N__10664\,
            I => \N__10617\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__10661\,
            I => \N__10617\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__10656\,
            I => \N__10617\
        );

    \I__2551\ : InMux
    port map (
            O => \N__10655\,
            I => \N__10612\
        );

    \I__2550\ : InMux
    port map (
            O => \N__10654\,
            I => \N__10612\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10607\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__10648\,
            I => \N__10607\
        );

    \I__2547\ : InMux
    port map (
            O => \N__10647\,
            I => \N__10604\
        );

    \I__2546\ : InMux
    port map (
            O => \N__10646\,
            I => \N__10599\
        );

    \I__2545\ : InMux
    port map (
            O => \N__10645\,
            I => \N__10599\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10596\
        );

    \I__2543\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10591\
        );

    \I__2542\ : InMux
    port map (
            O => \N__10640\,
            I => \N__10591\
        );

    \I__2541\ : InMux
    port map (
            O => \N__10639\,
            I => \N__10588\
        );

    \I__2540\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10585\
        );

    \I__2539\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10582\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__10626\,
            I => \N__10575\
        );

    \I__2537\ : Span4Mux_h
    port map (
            O => \N__10617\,
            I => \N__10575\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__10612\,
            I => \N__10575\
        );

    \I__2535\ : Span4Mux_v
    port map (
            O => \N__10607\,
            I => \N__10570\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__10604\,
            I => \N__10567\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__10599\,
            I => \N__10564\
        );

    \I__2532\ : Span4Mux_h
    port map (
            O => \N__10596\,
            I => \N__10555\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10555\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10588\,
            I => \N__10555\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10555\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10552\
        );

    \I__2527\ : Span4Mux_v
    port map (
            O => \N__10575\,
            I => \N__10549\
        );

    \I__2526\ : InMux
    port map (
            O => \N__10574\,
            I => \N__10546\
        );

    \I__2525\ : InMux
    port map (
            O => \N__10573\,
            I => \N__10543\
        );

    \I__2524\ : Span4Mux_h
    port map (
            O => \N__10570\,
            I => \N__10536\
        );

    \I__2523\ : Span4Mux_v
    port map (
            O => \N__10567\,
            I => \N__10536\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__10564\,
            I => \N__10536\
        );

    \I__2521\ : Span4Mux_h
    port map (
            O => \N__10555\,
            I => \N__10533\
        );

    \I__2520\ : Span4Mux_h
    port map (
            O => \N__10552\,
            I => \N__10528\
        );

    \I__2519\ : Span4Mux_h
    port map (
            O => \N__10549\,
            I => \N__10528\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10546\,
            I => \CPU_CYCLE\
        );

    \I__2517\ : LocalMux
    port map (
            O => \N__10543\,
            I => \CPU_CYCLE\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__10536\,
            I => \CPU_CYCLE\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__10533\,
            I => \CPU_CYCLE\
        );

    \I__2514\ : Odrv4
    port map (
            O => \N__10528\,
            I => \CPU_CYCLE\
        );

    \I__2513\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10513\
        );

    \I__2512\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10510\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__10513\,
            I => \N__10505\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10510\,
            I => \N__10505\
        );

    \I__2509\ : Span4Mux_v
    port map (
            O => \N__10505\,
            I => \N__10502\
        );

    \I__2508\ : Odrv4
    port map (
            O => \N__10502\,
            I => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\
        );

    \I__2507\ : CascadeMux
    port map (
            O => \N__10499\,
            I => \U712_BYTE_ENABLE.N_91_cascade_\
        );

    \I__2506\ : IoInMux
    port map (
            O => \N__10496\,
            I => \N__10493\
        );

    \I__2505\ : LocalMux
    port map (
            O => \N__10493\,
            I => \N__10490\
        );

    \I__2504\ : Span4Mux_s2_h
    port map (
            O => \N__10490\,
            I => \N__10487\
        );

    \I__2503\ : Sp12to4
    port map (
            O => \N__10487\,
            I => \N__10484\
        );

    \I__2502\ : Span12Mux_v
    port map (
            O => \N__10484\,
            I => \N__10481\
        );

    \I__2501\ : Span12Mux_h
    port map (
            O => \N__10481\,
            I => \N__10478\
        );

    \I__2500\ : Odrv12
    port map (
            O => \N__10478\,
            I => \N_51_i\
        );

    \I__2499\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10472\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__10472\,
            I => \U712_BYTE_ENABLE.N_89\
        );

    \I__2497\ : IoInMux
    port map (
            O => \N__10469\,
            I => \N__10466\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__10466\,
            I => \N__10463\
        );

    \I__2495\ : IoSpan4Mux
    port map (
            O => \N__10463\,
            I => \N__10460\
        );

    \I__2494\ : Span4Mux_s3_v
    port map (
            O => \N__10460\,
            I => \N__10457\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__10457\,
            I => \N_90_i\
        );

    \I__2492\ : IoInMux
    port map (
            O => \N__10454\,
            I => \N__10451\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10451\,
            I => \N__10448\
        );

    \I__2490\ : IoSpan4Mux
    port map (
            O => \N__10448\,
            I => \N__10445\
        );

    \I__2489\ : Span4Mux_s2_v
    port map (
            O => \N__10445\,
            I => \N__10442\
        );

    \I__2488\ : Span4Mux_v
    port map (
            O => \N__10442\,
            I => \N__10439\
        );

    \I__2487\ : Odrv4
    port map (
            O => \N__10439\,
            I => \N_92_i\
        );

    \I__2486\ : IoInMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10433\,
            I => \N__10430\
        );

    \I__2484\ : Span4Mux_s3_v
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__2483\ : Odrv4
    port map (
            O => \N__10427\,
            I => \N_91_i\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__10424\,
            I => \N__10420\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__10423\,
            I => \N__10417\
        );

    \I__2480\ : InMux
    port map (
            O => \N__10420\,
            I => \N__10413\
        );

    \I__2479\ : InMux
    port map (
            O => \N__10417\,
            I => \N__10408\
        );

    \I__2478\ : InMux
    port map (
            O => \N__10416\,
            I => \N__10408\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10413\,
            I => \N__10400\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__10408\,
            I => \N__10397\
        );

    \I__2475\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10394\
        );

    \I__2474\ : InMux
    port map (
            O => \N__10406\,
            I => \N__10385\
        );

    \I__2473\ : InMux
    port map (
            O => \N__10405\,
            I => \N__10385\
        );

    \I__2472\ : InMux
    port map (
            O => \N__10404\,
            I => \N__10385\
        );

    \I__2471\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10385\
        );

    \I__2470\ : Span4Mux_v
    port map (
            O => \N__10400\,
            I => \N__10382\
        );

    \I__2469\ : Sp12to4
    port map (
            O => \N__10397\,
            I => \N__10377\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__10394\,
            I => \N__10377\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10385\,
            I => \N__10374\
        );

    \I__2466\ : Span4Mux_v
    port map (
            O => \N__10382\,
            I => \N__10371\
        );

    \I__2465\ : Span12Mux_h
    port map (
            O => \N__10377\,
            I => \N__10368\
        );

    \I__2464\ : Span12Mux_v
    port map (
            O => \N__10374\,
            I => \N__10365\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10371\,
            I => \N__10362\
        );

    \I__2462\ : Span12Mux_v
    port map (
            O => \N__10368\,
            I => \N__10357\
        );

    \I__2461\ : Span12Mux_h
    port map (
            O => \N__10365\,
            I => \N__10357\
        );

    \I__2460\ : Sp12to4
    port map (
            O => \N__10362\,
            I => \N__10354\
        );

    \I__2459\ : Odrv12
    port map (
            O => \N__10357\,
            I => \SIZ_c_1\
        );

    \I__2458\ : Odrv12
    port map (
            O => \N__10354\,
            I => \SIZ_c_1\
        );

    \I__2457\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10342\
        );

    \I__2456\ : InMux
    port map (
            O => \N__10348\,
            I => \N__10342\
        );

    \I__2455\ : InMux
    port map (
            O => \N__10347\,
            I => \N__10339\
        );

    \I__2454\ : LocalMux
    port map (
            O => \N__10342\,
            I => \N__10332\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__10339\,
            I => \N__10329\
        );

    \I__2452\ : InMux
    port map (
            O => \N__10338\,
            I => \N__10320\
        );

    \I__2451\ : InMux
    port map (
            O => \N__10337\,
            I => \N__10320\
        );

    \I__2450\ : InMux
    port map (
            O => \N__10336\,
            I => \N__10320\
        );

    \I__2449\ : InMux
    port map (
            O => \N__10335\,
            I => \N__10320\
        );

    \I__2448\ : Span4Mux_v
    port map (
            O => \N__10332\,
            I => \N__10316\
        );

    \I__2447\ : Span4Mux_v
    port map (
            O => \N__10329\,
            I => \N__10313\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10320\,
            I => \N__10310\
        );

    \I__2445\ : InMux
    port map (
            O => \N__10319\,
            I => \N__10307\
        );

    \I__2444\ : Span4Mux_v
    port map (
            O => \N__10316\,
            I => \N__10300\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__10313\,
            I => \N__10300\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__10310\,
            I => \N__10300\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__10307\,
            I => \N__10297\
        );

    \I__2440\ : Sp12to4
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__2439\ : Sp12to4
    port map (
            O => \N__10297\,
            I => \N__10291\
        );

    \I__2438\ : Span12Mux_h
    port map (
            O => \N__10294\,
            I => \N__10286\
        );

    \I__2437\ : Span12Mux_v
    port map (
            O => \N__10291\,
            I => \N__10286\
        );

    \I__2436\ : Odrv12
    port map (
            O => \N__10286\,
            I => \A_c_1\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__10283\,
            I => \N__10278\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__10282\,
            I => \N__10273\
        );

    \I__2433\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10269\
        );

    \I__2432\ : InMux
    port map (
            O => \N__10278\,
            I => \N__10260\
        );

    \I__2431\ : InMux
    port map (
            O => \N__10277\,
            I => \N__10260\
        );

    \I__2430\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10260\
        );

    \I__2429\ : InMux
    port map (
            O => \N__10273\,
            I => \N__10260\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__10272\,
            I => \N__10255\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10269\,
            I => \N__10252\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10248\
        );

    \I__2425\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10245\
        );

    \I__2424\ : InMux
    port map (
            O => \N__10258\,
            I => \N__10239\
        );

    \I__2423\ : InMux
    port map (
            O => \N__10255\,
            I => \N__10239\
        );

    \I__2422\ : Span4Mux_v
    port map (
            O => \N__10252\,
            I => \N__10236\
        );

    \I__2421\ : InMux
    port map (
            O => \N__10251\,
            I => \N__10233\
        );

    \I__2420\ : Span4Mux_h
    port map (
            O => \N__10248\,
            I => \N__10230\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10227\
        );

    \I__2418\ : InMux
    port map (
            O => \N__10244\,
            I => \N__10224\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__10239\,
            I => \N__10217\
        );

    \I__2416\ : Sp12to4
    port map (
            O => \N__10236\,
            I => \N__10217\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__10233\,
            I => \N__10217\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__10230\,
            I => \N__10214\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__10227\,
            I => \N__10209\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10224\,
            I => \N__10209\
        );

    \I__2411\ : Span12Mux_h
    port map (
            O => \N__10217\,
            I => \N__10206\
        );

    \I__2410\ : Span4Mux_h
    port map (
            O => \N__10214\,
            I => \N__10203\
        );

    \I__2409\ : Sp12to4
    port map (
            O => \N__10209\,
            I => \N__10200\
        );

    \I__2408\ : Span12Mux_v
    port map (
            O => \N__10206\,
            I => \N__10197\
        );

    \I__2407\ : Sp12to4
    port map (
            O => \N__10203\,
            I => \N__10192\
        );

    \I__2406\ : Span12Mux_v
    port map (
            O => \N__10200\,
            I => \N__10192\
        );

    \I__2405\ : Odrv12
    port map (
            O => \N__10197\,
            I => \SIZ_c_0\
        );

    \I__2404\ : Odrv12
    port map (
            O => \N__10192\,
            I => \SIZ_c_0\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__10187\,
            I => \N__10182\
        );

    \I__2402\ : InMux
    port map (
            O => \N__10186\,
            I => \N__10174\
        );

    \I__2401\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10174\
        );

    \I__2400\ : InMux
    port map (
            O => \N__10182\,
            I => \N__10171\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__10181\,
            I => \N__10168\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__10180\,
            I => \N__10164\
        );

    \I__2397\ : CascadeMux
    port map (
            O => \N__10179\,
            I => \N__10161\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__10174\,
            I => \N__10157\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__10171\,
            I => \N__10154\
        );

    \I__2394\ : InMux
    port map (
            O => \N__10168\,
            I => \N__10151\
        );

    \I__2393\ : InMux
    port map (
            O => \N__10167\,
            I => \N__10142\
        );

    \I__2392\ : InMux
    port map (
            O => \N__10164\,
            I => \N__10142\
        );

    \I__2391\ : InMux
    port map (
            O => \N__10161\,
            I => \N__10142\
        );

    \I__2390\ : InMux
    port map (
            O => \N__10160\,
            I => \N__10142\
        );

    \I__2389\ : Span4Mux_h
    port map (
            O => \N__10157\,
            I => \N__10134\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__10154\,
            I => \N__10134\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__10151\,
            I => \N__10134\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__10142\,
            I => \N__10131\
        );

    \I__2385\ : InMux
    port map (
            O => \N__10141\,
            I => \N__10127\
        );

    \I__2384\ : Span4Mux_h
    port map (
            O => \N__10134\,
            I => \N__10124\
        );

    \I__2383\ : Span4Mux_v
    port map (
            O => \N__10131\,
            I => \N__10121\
        );

    \I__2382\ : InMux
    port map (
            O => \N__10130\,
            I => \N__10118\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__10127\,
            I => \N__10115\
        );

    \I__2380\ : Span4Mux_v
    port map (
            O => \N__10124\,
            I => \N__10112\
        );

    \I__2379\ : Sp12to4
    port map (
            O => \N__10121\,
            I => \N__10107\
        );

    \I__2378\ : LocalMux
    port map (
            O => \N__10118\,
            I => \N__10107\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10115\,
            I => \N__10104\
        );

    \I__2376\ : Sp12to4
    port map (
            O => \N__10112\,
            I => \N__10097\
        );

    \I__2375\ : Span12Mux_h
    port map (
            O => \N__10107\,
            I => \N__10097\
        );

    \I__2374\ : Sp12to4
    port map (
            O => \N__10104\,
            I => \N__10097\
        );

    \I__2373\ : Odrv12
    port map (
            O => \N__10097\,
            I => \A_c_0\
        );

    \I__2372\ : IoInMux
    port map (
            O => \N__10094\,
            I => \N__10091\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__10091\,
            I => \N__10088\
        );

    \I__2370\ : Span4Mux_s2_v
    port map (
            O => \N__10088\,
            I => \N__10085\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__10085\,
            I => \N__10082\
        );

    \I__2368\ : Span4Mux_v
    port map (
            O => \N__10082\,
            I => \N__10079\
        );

    \I__2367\ : Odrv4
    port map (
            O => \N__10079\,
            I => \N_89_i\
        );

    \I__2366\ : InMux
    port map (
            O => \N__10076\,
            I => \N__10072\
        );

    \I__2365\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10062\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__10069\,
            I => \N__10062\
        );

    \I__2362\ : InMux
    port map (
            O => \N__10068\,
            I => \N__10059\
        );

    \I__2361\ : InMux
    port map (
            O => \N__10067\,
            I => \N__10056\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__10062\,
            I => \N__10053\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__10059\,
            I => \N__10050\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__10056\,
            I => \N__10047\
        );

    \I__2357\ : Span4Mux_h
    port map (
            O => \N__10053\,
            I => \N__10042\
        );

    \I__2356\ : Span4Mux_v
    port map (
            O => \N__10050\,
            I => \N__10042\
        );

    \I__2355\ : Span12Mux_v
    port map (
            O => \N__10047\,
            I => \N__10039\
        );

    \I__2354\ : Span4Mux_v
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__2353\ : Span12Mux_h
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__2352\ : Sp12to4
    port map (
            O => \N__10036\,
            I => \N__10030\
        );

    \I__2351\ : Odrv12
    port map (
            O => \N__10033\,
            I => \DRA_c_3\
        );

    \I__2350\ : Odrv12
    port map (
            O => \N__10030\,
            I => \DRA_c_3\
        );

    \I__2349\ : InMux
    port map (
            O => \N__10025\,
            I => \N__10020\
        );

    \I__2348\ : InMux
    port map (
            O => \N__10024\,
            I => \N__10016\
        );

    \I__2347\ : InMux
    port map (
            O => \N__10023\,
            I => \N__10013\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__10020\,
            I => \N__10010\
        );

    \I__2345\ : InMux
    port map (
            O => \N__10019\,
            I => \N__10007\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__10016\,
            I => \N__10004\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__10013\,
            I => \N__10001\
        );

    \I__2342\ : Span4Mux_h
    port map (
            O => \N__10010\,
            I => \N__9996\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__10007\,
            I => \N__9996\
        );

    \I__2340\ : Span4Mux_v
    port map (
            O => \N__10004\,
            I => \N__9993\
        );

    \I__2339\ : Sp12to4
    port map (
            O => \N__10001\,
            I => \N__9988\
        );

    \I__2338\ : Sp12to4
    port map (
            O => \N__9996\,
            I => \N__9988\
        );

    \I__2337\ : Sp12to4
    port map (
            O => \N__9993\,
            I => \N__9985\
        );

    \I__2336\ : Span12Mux_v
    port map (
            O => \N__9988\,
            I => \N__9982\
        );

    \I__2335\ : Span12Mux_h
    port map (
            O => \N__9985\,
            I => \N__9979\
        );

    \I__2334\ : Span12Mux_h
    port map (
            O => \N__9982\,
            I => \N__9974\
        );

    \I__2333\ : Span12Mux_v
    port map (
            O => \N__9979\,
            I => \N__9974\
        );

    \I__2332\ : Odrv12
    port map (
            O => \N__9974\,
            I => \DRA_c_2\
        );

    \I__2331\ : InMux
    port map (
            O => \N__9971\,
            I => \N__9965\
        );

    \I__2330\ : InMux
    port map (
            O => \N__9970\,
            I => \N__9962\
        );

    \I__2329\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9956\
        );

    \I__2328\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9952\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9965\,
            I => \N__9945\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__9962\,
            I => \N__9942\
        );

    \I__2325\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9939\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9934\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9959\,
            I => \N__9934\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9956\,
            I => \N__9929\
        );

    \I__2321\ : InMux
    port map (
            O => \N__9955\,
            I => \N__9926\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__9952\,
            I => \N__9921\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9912\
        );

    \I__2318\ : InMux
    port map (
            O => \N__9950\,
            I => \N__9912\
        );

    \I__2317\ : InMux
    port map (
            O => \N__9949\,
            I => \N__9912\
        );

    \I__2316\ : InMux
    port map (
            O => \N__9948\,
            I => \N__9912\
        );

    \I__2315\ : Span4Mux_h
    port map (
            O => \N__9945\,
            I => \N__9904\
        );

    \I__2314\ : Span4Mux_h
    port map (
            O => \N__9942\,
            I => \N__9897\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__9939\,
            I => \N__9897\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__9934\,
            I => \N__9897\
        );

    \I__2311\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9892\
        );

    \I__2310\ : InMux
    port map (
            O => \N__9932\,
            I => \N__9892\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__9929\,
            I => \N__9889\
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__9926\,
            I => \N__9886\
        );

    \I__2307\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9881\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9881\
        );

    \I__2305\ : Span4Mux_h
    port map (
            O => \N__9921\,
            I => \N__9876\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9912\,
            I => \N__9876\
        );

    \I__2303\ : InMux
    port map (
            O => \N__9911\,
            I => \N__9867\
        );

    \I__2302\ : InMux
    port map (
            O => \N__9910\,
            I => \N__9867\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9909\,
            I => \N__9867\
        );

    \I__2300\ : InMux
    port map (
            O => \N__9908\,
            I => \N__9867\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9907\,
            I => \N__9864\
        );

    \I__2298\ : Span4Mux_h
    port map (
            O => \N__9904\,
            I => \N__9857\
        );

    \I__2297\ : Span4Mux_h
    port map (
            O => \N__9897\,
            I => \N__9857\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9892\,
            I => \N__9857\
        );

    \I__2295\ : Span4Mux_h
    port map (
            O => \N__9889\,
            I => \N__9854\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__9886\,
            I => \N__9851\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__9881\,
            I => \N__9848\
        );

    \I__2292\ : Sp12to4
    port map (
            O => \N__9876\,
            I => \N__9839\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__9867\,
            I => \N__9839\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9839\
        );

    \I__2289\ : Sp12to4
    port map (
            O => \N__9857\,
            I => \N__9839\
        );

    \I__2288\ : Sp12to4
    port map (
            O => \N__9854\,
            I => \N__9834\
        );

    \I__2287\ : Sp12to4
    port map (
            O => \N__9851\,
            I => \N__9834\
        );

    \I__2286\ : Span12Mux_h
    port map (
            O => \N__9848\,
            I => \N__9831\
        );

    \I__2285\ : Span12Mux_v
    port map (
            O => \N__9839\,
            I => \N__9828\
        );

    \I__2284\ : Span12Mux_h
    port map (
            O => \N__9834\,
            I => \N__9825\
        );

    \I__2283\ : Span12Mux_v
    port map (
            O => \N__9831\,
            I => \N__9820\
        );

    \I__2282\ : Span12Mux_h
    port map (
            O => \N__9828\,
            I => \N__9820\
        );

    \I__2281\ : Span12Mux_v
    port map (
            O => \N__9825\,
            I => \N__9817\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__9820\,
            I => \AGNUS_REV_c\
        );

    \I__2279\ : Odrv12
    port map (
            O => \N__9817\,
            I => \AGNUS_REV_c\
        );

    \I__2278\ : InMux
    port map (
            O => \N__9812\,
            I => \N__9809\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9806\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__9806\,
            I => \N__9803\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__9803\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\
        );

    \I__2274\ : ClkMux
    port map (
            O => \N__9800\,
            I => \N__9785\
        );

    \I__2273\ : ClkMux
    port map (
            O => \N__9799\,
            I => \N__9785\
        );

    \I__2272\ : ClkMux
    port map (
            O => \N__9798\,
            I => \N__9785\
        );

    \I__2271\ : ClkMux
    port map (
            O => \N__9797\,
            I => \N__9785\
        );

    \I__2270\ : ClkMux
    port map (
            O => \N__9796\,
            I => \N__9785\
        );

    \I__2269\ : GlobalMux
    port map (
            O => \N__9785\,
            I => \N__9782\
        );

    \I__2268\ : gio2CtrlBuf
    port map (
            O => \N__9782\,
            I => \C3_c_g\
        );

    \I__2267\ : CEMux
    port map (
            O => \N__9779\,
            I => \N__9749\
        );

    \I__2266\ : CEMux
    port map (
            O => \N__9778\,
            I => \N__9749\
        );

    \I__2265\ : CEMux
    port map (
            O => \N__9777\,
            I => \N__9749\
        );

    \I__2264\ : CEMux
    port map (
            O => \N__9776\,
            I => \N__9749\
        );

    \I__2263\ : CEMux
    port map (
            O => \N__9775\,
            I => \N__9749\
        );

    \I__2262\ : CEMux
    port map (
            O => \N__9774\,
            I => \N__9749\
        );

    \I__2261\ : CEMux
    port map (
            O => \N__9773\,
            I => \N__9749\
        );

    \I__2260\ : CEMux
    port map (
            O => \N__9772\,
            I => \N__9749\
        );

    \I__2259\ : CEMux
    port map (
            O => \N__9771\,
            I => \N__9749\
        );

    \I__2258\ : CEMux
    port map (
            O => \N__9770\,
            I => \N__9749\
        );

    \I__2257\ : GlobalMux
    port map (
            O => \N__9749\,
            I => \N__9746\
        );

    \I__2256\ : gio2CtrlBuf
    port map (
            O => \N__9746\,
            I => \DBRn_c_i_0_g\
        );

    \I__2255\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9740\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9720\
        );

    \I__2253\ : ClkMux
    port map (
            O => \N__9739\,
            I => \N__9662\
        );

    \I__2252\ : ClkMux
    port map (
            O => \N__9738\,
            I => \N__9662\
        );

    \I__2251\ : ClkMux
    port map (
            O => \N__9737\,
            I => \N__9662\
        );

    \I__2250\ : ClkMux
    port map (
            O => \N__9736\,
            I => \N__9662\
        );

    \I__2249\ : ClkMux
    port map (
            O => \N__9735\,
            I => \N__9662\
        );

    \I__2248\ : ClkMux
    port map (
            O => \N__9734\,
            I => \N__9662\
        );

    \I__2247\ : ClkMux
    port map (
            O => \N__9733\,
            I => \N__9662\
        );

    \I__2246\ : ClkMux
    port map (
            O => \N__9732\,
            I => \N__9662\
        );

    \I__2245\ : ClkMux
    port map (
            O => \N__9731\,
            I => \N__9662\
        );

    \I__2244\ : ClkMux
    port map (
            O => \N__9730\,
            I => \N__9662\
        );

    \I__2243\ : ClkMux
    port map (
            O => \N__9729\,
            I => \N__9662\
        );

    \I__2242\ : ClkMux
    port map (
            O => \N__9728\,
            I => \N__9662\
        );

    \I__2241\ : ClkMux
    port map (
            O => \N__9727\,
            I => \N__9662\
        );

    \I__2240\ : ClkMux
    port map (
            O => \N__9726\,
            I => \N__9662\
        );

    \I__2239\ : ClkMux
    port map (
            O => \N__9725\,
            I => \N__9662\
        );

    \I__2238\ : ClkMux
    port map (
            O => \N__9724\,
            I => \N__9662\
        );

    \I__2237\ : ClkMux
    port map (
            O => \N__9723\,
            I => \N__9662\
        );

    \I__2236\ : Glb2LocalMux
    port map (
            O => \N__9720\,
            I => \N__9662\
        );

    \I__2235\ : ClkMux
    port map (
            O => \N__9719\,
            I => \N__9662\
        );

    \I__2234\ : ClkMux
    port map (
            O => \N__9718\,
            I => \N__9662\
        );

    \I__2233\ : ClkMux
    port map (
            O => \N__9717\,
            I => \N__9662\
        );

    \I__2232\ : ClkMux
    port map (
            O => \N__9716\,
            I => \N__9662\
        );

    \I__2231\ : ClkMux
    port map (
            O => \N__9715\,
            I => \N__9662\
        );

    \I__2230\ : ClkMux
    port map (
            O => \N__9714\,
            I => \N__9662\
        );

    \I__2229\ : ClkMux
    port map (
            O => \N__9713\,
            I => \N__9662\
        );

    \I__2228\ : GlobalMux
    port map (
            O => \N__9662\,
            I => \CLK80_PLL\
        );

    \I__2227\ : CEMux
    port map (
            O => \N__9659\,
            I => \N__9656\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__9656\,
            I => \N__9651\
        );

    \I__2225\ : CEMux
    port map (
            O => \N__9655\,
            I => \N__9648\
        );

    \I__2224\ : CEMux
    port map (
            O => \N__9654\,
            I => \N__9644\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__9651\,
            I => \N__9639\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9648\,
            I => \N__9639\
        );

    \I__2221\ : CEMux
    port map (
            O => \N__9647\,
            I => \N__9636\
        );

    \I__2220\ : LocalMux
    port map (
            O => \N__9644\,
            I => \N__9631\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__9639\,
            I => \N__9631\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__9636\,
            I => \N__9628\
        );

    \I__2217\ : Odrv4
    port map (
            O => \N__9631\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__9628\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_0\
        );

    \I__2215\ : InMux
    port map (
            O => \N__9623\,
            I => \N__9620\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__9620\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\
        );

    \I__2213\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9614\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9614\,
            I => \N__9608\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9603\
        );

    \I__2210\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9603\
        );

    \I__2209\ : InMux
    port map (
            O => \N__9611\,
            I => \N__9600\
        );

    \I__2208\ : Span4Mux_v
    port map (
            O => \N__9608\,
            I => \N__9597\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__9603\,
            I => \N__9592\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__9600\,
            I => \N__9592\
        );

    \I__2205\ : Span4Mux_v
    port map (
            O => \N__9597\,
            I => \N__9589\
        );

    \I__2204\ : Sp12to4
    port map (
            O => \N__9592\,
            I => \N__9586\
        );

    \I__2203\ : Sp12to4
    port map (
            O => \N__9589\,
            I => \N__9583\
        );

    \I__2202\ : Span12Mux_v
    port map (
            O => \N__9586\,
            I => \N__9580\
        );

    \I__2201\ : Span12Mux_h
    port map (
            O => \N__9583\,
            I => \N__9577\
        );

    \I__2200\ : Span12Mux_h
    port map (
            O => \N__9580\,
            I => \N__9574\
        );

    \I__2199\ : Odrv12
    port map (
            O => \N__9577\,
            I => \DRA_c_5\
        );

    \I__2198\ : Odrv12
    port map (
            O => \N__9574\,
            I => \DRA_c_5\
        );

    \I__2197\ : InMux
    port map (
            O => \N__9569\,
            I => \N__9563\
        );

    \I__2196\ : InMux
    port map (
            O => \N__9568\,
            I => \N__9563\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__9563\,
            I => \N__9560\
        );

    \I__2194\ : Span4Mux_h
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__2193\ : Odrv4
    port map (
            O => \N__9557\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\
        );

    \I__2192\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9550\
        );

    \I__2191\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9547\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__9550\,
            I => \N__9541\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__9547\,
            I => \N__9541\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9546\,
            I => \N__9538\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__9541\,
            I => \N__9532\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__9538\,
            I => \N__9532\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9529\
        );

    \I__2184\ : Span4Mux_v
    port map (
            O => \N__9532\,
            I => \N__9526\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__9529\,
            I => \N__9523\
        );

    \I__2182\ : Span4Mux_v
    port map (
            O => \N__9526\,
            I => \N__9520\
        );

    \I__2181\ : Span12Mux_v
    port map (
            O => \N__9523\,
            I => \N__9517\
        );

    \I__2180\ : Sp12to4
    port map (
            O => \N__9520\,
            I => \N__9514\
        );

    \I__2179\ : Span12Mux_h
    port map (
            O => \N__9517\,
            I => \N__9511\
        );

    \I__2178\ : Span12Mux_h
    port map (
            O => \N__9514\,
            I => \N__9508\
        );

    \I__2177\ : Odrv12
    port map (
            O => \N__9511\,
            I => \DRA_c_4\
        );

    \I__2176\ : Odrv12
    port map (
            O => \N__9508\,
            I => \DRA_c_4\
        );

    \I__2175\ : InMux
    port map (
            O => \N__9503\,
            I => \N__9500\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9500\,
            I => \N__9497\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__9497\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\
        );

    \I__2172\ : InMux
    port map (
            O => \N__9494\,
            I => \N__9491\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__9491\,
            I => \N__9488\
        );

    \I__2170\ : Odrv4
    port map (
            O => \N__9488\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\
        );

    \I__2169\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9481\
        );

    \I__2168\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9478\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__9481\,
            I => \N__9473\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9470\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9477\,
            I => \N__9465\
        );

    \I__2164\ : InMux
    port map (
            O => \N__9476\,
            I => \N__9465\
        );

    \I__2163\ : Span4Mux_v
    port map (
            O => \N__9473\,
            I => \N__9462\
        );

    \I__2162\ : Span4Mux_v
    port map (
            O => \N__9470\,
            I => \N__9459\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9456\
        );

    \I__2160\ : Sp12to4
    port map (
            O => \N__9462\,
            I => \N__9451\
        );

    \I__2159\ : Sp12to4
    port map (
            O => \N__9459\,
            I => \N__9451\
        );

    \I__2158\ : Span12Mux_v
    port map (
            O => \N__9456\,
            I => \N__9448\
        );

    \I__2157\ : Span12Mux_h
    port map (
            O => \N__9451\,
            I => \N__9445\
        );

    \I__2156\ : Span12Mux_h
    port map (
            O => \N__9448\,
            I => \N__9442\
        );

    \I__2155\ : Odrv12
    port map (
            O => \N__9445\,
            I => \DRA_c_8\
        );

    \I__2154\ : Odrv12
    port map (
            O => \N__9442\,
            I => \DRA_c_8\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__9437\,
            I => \N__9434\
        );

    \I__2152\ : InMux
    port map (
            O => \N__9434\,
            I => \N__9431\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__9431\,
            I => \N__9428\
        );

    \I__2150\ : Odrv4
    port map (
            O => \N__9428\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\
        );

    \I__2149\ : InMux
    port map (
            O => \N__9425\,
            I => \N__9422\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2147\ : Span12Mux_h
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__2146\ : Odrv12
    port map (
            O => \N__9416\,
            I => \RAS0n_c\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__9413\,
            I => \N__9410\
        );

    \I__2144\ : InMux
    port map (
            O => \N__9410\,
            I => \N__9407\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9407\,
            I => \N__9403\
        );

    \I__2142\ : InMux
    port map (
            O => \N__9406\,
            I => \N__9400\
        );

    \I__2141\ : Span4Mux_v
    port map (
            O => \N__9403\,
            I => \N__9393\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__9400\,
            I => \N__9393\
        );

    \I__2139\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9388\
        );

    \I__2138\ : InMux
    port map (
            O => \N__9398\,
            I => \N__9388\
        );

    \I__2137\ : Span4Mux_h
    port map (
            O => \N__9393\,
            I => \N__9383\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__9388\,
            I => \N__9383\
        );

    \I__2135\ : Span4Mux_h
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__2133\ : Sp12to4
    port map (
            O => \N__9377\,
            I => \N__9374\
        );

    \I__2132\ : Span12Mux_v
    port map (
            O => \N__9374\,
            I => \N__9371\
        );

    \I__2131\ : Odrv12
    port map (
            O => \N__9371\,
            I => \DRA_c_9\
        );

    \I__2130\ : InMux
    port map (
            O => \N__9368\,
            I => \N__9365\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__9365\,
            I => \N__9362\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__9362\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\
        );

    \I__2127\ : InMux
    port map (
            O => \N__9359\,
            I => \N__9352\
        );

    \I__2126\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__2125\ : InMux
    port map (
            O => \N__9357\,
            I => \N__9348\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__9352\,
            I => \N__9345\
        );

    \I__2123\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9342\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__9348\,
            I => \N__9335\
        );

    \I__2121\ : Sp12to4
    port map (
            O => \N__9345\,
            I => \N__9335\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__9342\,
            I => \N__9335\
        );

    \I__2119\ : Span12Mux_v
    port map (
            O => \N__9335\,
            I => \N__9332\
        );

    \I__2118\ : Span12Mux_h
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__2117\ : Odrv12
    port map (
            O => \N__9329\,
            I => \DRA_c_6\
        );

    \I__2116\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9318\
        );

    \I__2115\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9318\
        );

    \I__2114\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9315\
        );

    \I__2113\ : InMux
    port map (
            O => \N__9323\,
            I => \N__9312\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__9318\,
            I => \N__9309\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__9315\,
            I => \N__9304\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9304\
        );

    \I__2109\ : Span4Mux_v
    port map (
            O => \N__9309\,
            I => \N__9301\
        );

    \I__2108\ : Span4Mux_v
    port map (
            O => \N__9304\,
            I => \N__9298\
        );

    \I__2107\ : Sp12to4
    port map (
            O => \N__9301\,
            I => \N__9295\
        );

    \I__2106\ : Sp12to4
    port map (
            O => \N__9298\,
            I => \N__9292\
        );

    \I__2105\ : Span12Mux_h
    port map (
            O => \N__9295\,
            I => \N__9289\
        );

    \I__2104\ : Span12Mux_h
    port map (
            O => \N__9292\,
            I => \N__9286\
        );

    \I__2103\ : Odrv12
    port map (
            O => \N__9289\,
            I => \DRA_c_7\
        );

    \I__2102\ : Odrv12
    port map (
            O => \N__9286\,
            I => \DRA_c_7\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__9281\,
            I => \N__9278\
        );

    \I__2100\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__9275\,
            I => \N__9272\
        );

    \I__2098\ : Odrv12
    port map (
            O => \N__9272\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\
        );

    \I__2097\ : IoInMux
    port map (
            O => \N__9269\,
            I => \N__9266\
        );

    \I__2096\ : LocalMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__2095\ : Span4Mux_s2_h
    port map (
            O => \N__9263\,
            I => \N__9260\
        );

    \I__2094\ : Sp12to4
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__2093\ : Span12Mux_v
    port map (
            O => \N__9257\,
            I => \N__9254\
        );

    \I__2092\ : Span12Mux_v
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__2091\ : Span12Mux_h
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__2090\ : Odrv12
    port map (
            O => \N__9248\,
            I => \N_50_i\
        );

    \I__2089\ : IoInMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__9242\,
            I => \N__9239\
        );

    \I__2087\ : IoSpan4Mux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__2086\ : Sp12to4
    port map (
            O => \N__9236\,
            I => \N__9233\
        );

    \I__2085\ : Span12Mux_s7_v
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__2084\ : Odrv12
    port map (
            O => \N__9230\,
            I => \WEn_c\
        );

    \I__2083\ : IoInMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9221\
        );

    \I__2081\ : Span4Mux_s3_v
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__2080\ : Span4Mux_v
    port map (
            O => \N__9218\,
            I => \N__9215\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__2078\ : Odrv4
    port map (
            O => \N__9212\,
            I => \RASn_c\
        );

    \I__2077\ : IoInMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__9206\,
            I => \N__9203\
        );

    \I__2075\ : Span4Mux_s0_v
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__2074\ : Sp12to4
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__2073\ : Span12Mux_h
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__2072\ : Odrv12
    port map (
            O => \N__9194\,
            I => \CRCSn_c\
        );

    \I__2071\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9187\
        );

    \I__2070\ : InMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__9187\,
            I => \N__9180\
        );

    \I__2068\ : LocalMux
    port map (
            O => \N__9184\,
            I => \N__9177\
        );

    \I__2067\ : InMux
    port map (
            O => \N__9183\,
            I => \N__9174\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__9180\,
            I => \N__9164\
        );

    \I__2065\ : Span4Mux_h
    port map (
            O => \N__9177\,
            I => \N__9164\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9164\
        );

    \I__2063\ : InMux
    port map (
            O => \N__9173\,
            I => \N__9161\
        );

    \I__2062\ : InMux
    port map (
            O => \N__9172\,
            I => \N__9158\
        );

    \I__2061\ : InMux
    port map (
            O => \N__9171\,
            I => \N__9155\
        );

    \I__2060\ : Span4Mux_h
    port map (
            O => \N__9164\,
            I => \N__9152\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__9161\,
            I => \N__9149\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9158\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__9155\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__9152\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2055\ : Odrv12
    port map (
            O => \N__9149\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__9140\,
            I => \N__9131\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__9139\,
            I => \N__9128\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__9138\,
            I => \N__9125\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__9137\,
            I => \N__9119\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__9136\,
            I => \N__9113\
        );

    \I__2049\ : InMux
    port map (
            O => \N__9135\,
            I => \N__9110\
        );

    \I__2048\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9107\
        );

    \I__2047\ : InMux
    port map (
            O => \N__9131\,
            I => \N__9104\
        );

    \I__2046\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9097\
        );

    \I__2045\ : InMux
    port map (
            O => \N__9125\,
            I => \N__9097\
        );

    \I__2044\ : InMux
    port map (
            O => \N__9124\,
            I => \N__9097\
        );

    \I__2043\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9094\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__9122\,
            I => \N__9091\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9119\,
            I => \N__9087\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9118\,
            I => \N__9080\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9117\,
            I => \N__9080\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9116\,
            I => \N__9080\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9077\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9110\,
            I => \N__9072\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__9107\,
            I => \N__9069\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9059\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9097\,
            I => \N__9059\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9094\,
            I => \N__9059\
        );

    \I__2031\ : InMux
    port map (
            O => \N__9091\,
            I => \N__9054\
        );

    \I__2030\ : InMux
    port map (
            O => \N__9090\,
            I => \N__9054\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9087\,
            I => \N__9047\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__9080\,
            I => \N__9047\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__9077\,
            I => \N__9047\
        );

    \I__2026\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9044\
        );

    \I__2025\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9041\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__9072\,
            I => \N__9032\
        );

    \I__2023\ : Span4Mux_h
    port map (
            O => \N__9069\,
            I => \N__9032\
        );

    \I__2022\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9025\
        );

    \I__2021\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9025\
        );

    \I__2020\ : InMux
    port map (
            O => \N__9066\,
            I => \N__9025\
        );

    \I__2019\ : Span4Mux_v
    port map (
            O => \N__9059\,
            I => \N__9020\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9020\
        );

    \I__2017\ : Span4Mux_v
    port map (
            O => \N__9047\,
            I => \N__9017\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__9044\,
            I => \N__9014\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__9041\,
            I => \N__9011\
        );

    \I__2014\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9002\
        );

    \I__2013\ : InMux
    port map (
            O => \N__9039\,
            I => \N__9002\
        );

    \I__2012\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9002\
        );

    \I__2011\ : InMux
    port map (
            O => \N__9037\,
            I => \N__9002\
        );

    \I__2010\ : Span4Mux_h
    port map (
            O => \N__9032\,
            I => \N__8997\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__9025\,
            I => \N__8997\
        );

    \I__2008\ : Span4Mux_h
    port map (
            O => \N__9020\,
            I => \N__8994\
        );

    \I__2007\ : Odrv4
    port map (
            O => \N__9017\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2006\ : Odrv4
    port map (
            O => \N__9014\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__9011\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__9002\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2003\ : Odrv4
    port map (
            O => \N__8997\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__8994\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\
        );

    \I__2001\ : CascadeMux
    port map (
            O => \N__8981\,
            I => \N__8976\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__8980\,
            I => \N__8973\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8979\,
            I => \N__8969\
        );

    \I__1998\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8966\
        );

    \I__1997\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8963\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__8972\,
            I => \N__8960\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__8969\,
            I => \N__8955\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8955\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8963\,
            I => \N__8952\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8960\,
            I => \N__8949\
        );

    \I__1991\ : Span4Mux_v
    port map (
            O => \N__8955\,
            I => \N__8946\
        );

    \I__1990\ : Span4Mux_v
    port map (
            O => \N__8952\,
            I => \N__8941\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8949\,
            I => \N__8941\
        );

    \I__1988\ : Odrv4
    port map (
            O => \N__8946\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__8941\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\
        );

    \I__1986\ : InMux
    port map (
            O => \N__8936\,
            I => \N__8932\
        );

    \I__1985\ : InMux
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8932\,
            I => \N__8923\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8923\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8928\,
            I => \N__8920\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__8923\,
            I => \N__8916\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8911\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8908\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__8916\,
            I => \N__8905\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8915\,
            I => \N__8902\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8914\,
            I => \N__8899\
        );

    \I__1975\ : Span4Mux_v
    port map (
            O => \N__8911\,
            I => \N__8894\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__8908\,
            I => \N__8894\
        );

    \I__1973\ : Odrv4
    port map (
            O => \N__8905\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__8902\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__8899\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__8894\,
            I => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\
        );

    \I__1969\ : IoInMux
    port map (
            O => \N__8885\,
            I => \N__8882\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8882\,
            I => \N__8879\
        );

    \I__1967\ : Span12Mux_s10_v
    port map (
            O => \N__8879\,
            I => \N__8876\
        );

    \I__1966\ : Odrv12
    port map (
            O => \N__8876\,
            I => \CMA_c_10\
        );

    \I__1965\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8870\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8870\,
            I => \N__8867\
        );

    \I__1963\ : Span4Mux_v
    port map (
            O => \N__8867\,
            I => \N__8864\
        );

    \I__1962\ : Span4Mux_v
    port map (
            O => \N__8864\,
            I => \N__8861\
        );

    \I__1961\ : Sp12to4
    port map (
            O => \N__8861\,
            I => \N__8858\
        );

    \I__1960\ : Span12Mux_h
    port map (
            O => \N__8858\,
            I => \N__8855\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__8855\,
            I => \A_c_17\
        );

    \I__1958\ : IoInMux
    port map (
            O => \N__8852\,
            I => \N__8849\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8846\
        );

    \I__1956\ : IoSpan4Mux
    port map (
            O => \N__8846\,
            I => \N__8843\
        );

    \I__1955\ : IoSpan4Mux
    port map (
            O => \N__8843\,
            I => \N__8840\
        );

    \I__1954\ : Span4Mux_s3_h
    port map (
            O => \N__8840\,
            I => \N__8837\
        );

    \I__1953\ : Sp12to4
    port map (
            O => \N__8837\,
            I => \N__8834\
        );

    \I__1952\ : Odrv12
    port map (
            O => \N__8834\,
            I => \CMA_c_8\
        );

    \I__1951\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8828\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8825\
        );

    \I__1949\ : Odrv12
    port map (
            O => \N__8825\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\
        );

    \I__1948\ : IoInMux
    port map (
            O => \N__8822\,
            I => \N__8819\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__8819\,
            I => \N__8816\
        );

    \I__1946\ : Span12Mux_s2_h
    port map (
            O => \N__8816\,
            I => \N__8813\
        );

    \I__1945\ : Span12Mux_h
    port map (
            O => \N__8813\,
            I => \N__8810\
        );

    \I__1944\ : Odrv12
    port map (
            O => \N__8810\,
            I => \CMA_c_3\
        );

    \I__1943\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8804\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__8804\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\
        );

    \I__1941\ : IoInMux
    port map (
            O => \N__8801\,
            I => \N__8798\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8798\,
            I => \N__8795\
        );

    \I__1939\ : Span4Mux_s2_h
    port map (
            O => \N__8795\,
            I => \N__8792\
        );

    \I__1938\ : Sp12to4
    port map (
            O => \N__8792\,
            I => \N__8789\
        );

    \I__1937\ : Span12Mux_s10_v
    port map (
            O => \N__8789\,
            I => \N__8786\
        );

    \I__1936\ : Span12Mux_h
    port map (
            O => \N__8786\,
            I => \N__8783\
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__8783\,
            I => \CMA_c_6\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8780\,
            I => \N__8770\
        );

    \I__1933\ : InMux
    port map (
            O => \N__8779\,
            I => \N__8765\
        );

    \I__1932\ : InMux
    port map (
            O => \N__8778\,
            I => \N__8765\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8777\,
            I => \N__8762\
        );

    \I__1930\ : InMux
    port map (
            O => \N__8776\,
            I => \N__8757\
        );

    \I__1929\ : InMux
    port map (
            O => \N__8775\,
            I => \N__8757\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__8774\,
            I => \N__8754\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__8773\,
            I => \N__8751\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8770\,
            I => \N__8741\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8765\,
            I => \N__8741\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8741\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__8757\,
            I => \N__8741\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8734\
        );

    \I__1921\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8734\
        );

    \I__1920\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8734\
        );

    \I__1919\ : Odrv12
    port map (
            O => \N__8741\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__8734\,
            I => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__8729\,
            I => \N__8722\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__8728\,
            I => \N__8719\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__8727\,
            I => \N__8715\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__8726\,
            I => \N__8712\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8725\,
            I => \N__8705\
        );

    \I__1912\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8705\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8719\,
            I => \N__8705\
        );

    \I__1910\ : InMux
    port map (
            O => \N__8718\,
            I => \N__8698\
        );

    \I__1909\ : InMux
    port map (
            O => \N__8715\,
            I => \N__8698\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8698\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__8705\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__8698\,
            I => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\
        );

    \I__1905\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__8690\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\
        );

    \I__1903\ : IoInMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__8684\,
            I => \N__8681\
        );

    \I__1901\ : IoSpan4Mux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__1900\ : Span4Mux_s3_h
    port map (
            O => \N__8678\,
            I => \N__8675\
        );

    \I__1899\ : Sp12to4
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1898\ : Span12Mux_h
    port map (
            O => \N__8672\,
            I => \N__8669\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__8669\,
            I => \CMA_c_4\
        );

    \I__1896\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__8660\,
            I => \N__8657\
        );

    \I__1893\ : Span4Mux_v
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__1892\ : Sp12to4
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__1891\ : Span12Mux_h
    port map (
            O => \N__8651\,
            I => \N__8648\
        );

    \I__1890\ : Odrv12
    port map (
            O => \N__8648\,
            I => \A_c_19\
        );

    \I__1889\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8642\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8638\
        );

    \I__1887\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8635\
        );

    \I__1886\ : Span4Mux_v
    port map (
            O => \N__8638\,
            I => \N__8630\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__8635\,
            I => \N__8627\
        );

    \I__1884\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8622\
        );

    \I__1883\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8622\
        );

    \I__1882\ : Odrv4
    port map (
            O => \N__8630\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1881\ : Odrv12
    port map (
            O => \N__8627\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__8622\,
            I => \U712_CHIP_RAM.CMA_5_0_8\
        );

    \I__1879\ : IoInMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__8612\,
            I => \N__8609\
        );

    \I__1877\ : IoSpan4Mux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__1876\ : IoSpan4Mux
    port map (
            O => \N__8606\,
            I => \N__8603\
        );

    \I__1875\ : Span4Mux_s3_h
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__1874\ : Sp12to4
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__1873\ : Odrv12
    port map (
            O => \N__8597\,
            I => \CMA_c_9\
        );

    \I__1872\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__8591\,
            I => \N__8588\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__8588\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\
        );

    \I__1869\ : InMux
    port map (
            O => \N__8585\,
            I => \N__8579\
        );

    \I__1868\ : InMux
    port map (
            O => \N__8584\,
            I => \N__8579\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__8579\,
            I => \N__8576\
        );

    \I__1866\ : Odrv4
    port map (
            O => \N__8576\,
            I => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\
        );

    \I__1865\ : InMux
    port map (
            O => \N__8573\,
            I => \N__8570\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__1863\ : Odrv4
    port map (
            O => \N__8567\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\
        );

    \I__1862\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8558\
        );

    \I__1861\ : InMux
    port map (
            O => \N__8563\,
            I => \N__8558\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8553\
        );

    \I__1859\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8548\
        );

    \I__1858\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8548\
        );

    \I__1857\ : Span4Mux_v
    port map (
            O => \N__8553\,
            I => \N__8545\
        );

    \I__1856\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8542\
        );

    \I__1855\ : Span4Mux_h
    port map (
            O => \N__8545\,
            I => \N__8539\
        );

    \I__1854\ : Span12Mux_h
    port map (
            O => \N__8542\,
            I => \N__8534\
        );

    \I__1853\ : Sp12to4
    port map (
            O => \N__8539\,
            I => \N__8534\
        );

    \I__1852\ : Span12Mux_v
    port map (
            O => \N__8534\,
            I => \N__8531\
        );

    \I__1851\ : Odrv12
    port map (
            O => \N__8531\,
            I => \DRA_c_1\
        );

    \I__1850\ : InMux
    port map (
            O => \N__8528\,
            I => \N__8525\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__8522\,
            I => \N__8518\
        );

    \I__1847\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1846\ : Sp12to4
    port map (
            O => \N__8518\,
            I => \N__8510\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__8515\,
            I => \N__8510\
        );

    \I__1844\ : Span12Mux_h
    port map (
            O => \N__8510\,
            I => \N__8507\
        );

    \I__1843\ : Span12Mux_v
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__1842\ : Odrv12
    port map (
            O => \N__8504\,
            I => \DRA_c_0\
        );

    \I__1841\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__8498\,
            I => \N__8495\
        );

    \I__1839\ : Odrv12
    port map (
            O => \N__8495\,
            I => \U712_CHIP_RAM.DMA_AZ0Z1\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__8492\,
            I => \N__8485\
        );

    \I__1837\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8481\
        );

    \I__1836\ : InMux
    port map (
            O => \N__8490\,
            I => \N__8476\
        );

    \I__1835\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8469\
        );

    \I__1834\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8469\
        );

    \I__1833\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8469\
        );

    \I__1832\ : InMux
    port map (
            O => \N__8484\,
            I => \N__8466\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__8481\,
            I => \N__8463\
        );

    \I__1830\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8458\
        );

    \I__1829\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8458\
        );

    \I__1828\ : LocalMux
    port map (
            O => \N__8476\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__8469\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__8466\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1825\ : Odrv4
    port map (
            O => \N__8463\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__8458\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_0\
        );

    \I__1823\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8444\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__8444\,
            I => \U712_REG_SM.N_369\
        );

    \I__1821\ : IoInMux
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__1819\ : IoSpan4Mux
    port map (
            O => \N__8435\,
            I => \N__8432\
        );

    \I__1818\ : Span4Mux_s3_v
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__1817\ : Sp12to4
    port map (
            O => \N__8429\,
            I => \N__8425\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__1815\ : Span12Mux_h
    port map (
            O => \N__8425\,
            I => \N__8417\
        );

    \I__1814\ : InMux
    port map (
            O => \N__8422\,
            I => \N__8414\
        );

    \I__1813\ : InMux
    port map (
            O => \N__8421\,
            I => \N__8411\
        );

    \I__1812\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8408\
        );

    \I__1811\ : Odrv12
    port map (
            O => \N__8417\,
            I => \UDSn_c\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__8414\,
            I => \UDSn_c\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__8411\,
            I => \UDSn_c\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__8408\,
            I => \UDSn_c\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8399\,
            I => \N__8395\
        );

    \I__1806\ : InMux
    port map (
            O => \N__8398\,
            I => \N__8385\
        );

    \I__1805\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8385\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8394\,
            I => \N__8385\
        );

    \I__1803\ : InMux
    port map (
            O => \N__8393\,
            I => \N__8382\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__8392\,
            I => \N__8379\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__8385\,
            I => \N__8370\
        );

    \I__1800\ : LocalMux
    port map (
            O => \N__8382\,
            I => \N__8370\
        );

    \I__1799\ : InMux
    port map (
            O => \N__8379\,
            I => \N__8367\
        );

    \I__1798\ : InMux
    port map (
            O => \N__8378\,
            I => \N__8364\
        );

    \I__1797\ : InMux
    port map (
            O => \N__8377\,
            I => \N__8359\
        );

    \I__1796\ : InMux
    port map (
            O => \N__8376\,
            I => \N__8359\
        );

    \I__1795\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8356\
        );

    \I__1794\ : Span4Mux_h
    port map (
            O => \N__8370\,
            I => \N__8353\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__8367\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__8364\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8359\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__8356\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__8353\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_2\
        );

    \I__1788\ : InMux
    port map (
            O => \N__8342\,
            I => \N__8339\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__8339\,
            I => \U712_REG_SM.N_465\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__8336\,
            I => \N__8333\
        );

    \I__1785\ : InMux
    port map (
            O => \N__8333\,
            I => \N__8328\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__8332\,
            I => \N__8323\
        );

    \I__1783\ : InMux
    port map (
            O => \N__8331\,
            I => \N__8320\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__8328\,
            I => \N__8314\
        );

    \I__1781\ : InMux
    port map (
            O => \N__8327\,
            I => \N__8309\
        );

    \I__1780\ : InMux
    port map (
            O => \N__8326\,
            I => \N__8309\
        );

    \I__1779\ : InMux
    port map (
            O => \N__8323\,
            I => \N__8306\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__8320\,
            I => \N__8303\
        );

    \I__1777\ : InMux
    port map (
            O => \N__8319\,
            I => \N__8300\
        );

    \I__1776\ : InMux
    port map (
            O => \N__8318\,
            I => \N__8295\
        );

    \I__1775\ : InMux
    port map (
            O => \N__8317\,
            I => \N__8295\
        );

    \I__1774\ : Odrv4
    port map (
            O => \N__8314\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__8309\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__8306\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__8303\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__8300\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__8295\,
            I => \U712_REG_SM.C1_SYNCZ0Z_1\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__8282\,
            I => \N__8277\
        );

    \I__1767\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8274\
        );

    \I__1766\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8271\
        );

    \I__1765\ : InMux
    port map (
            O => \N__8277\,
            I => \N__8268\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__8274\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__8271\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__8268\,
            I => \U712_REG_SM.REG_CYCLE_STARTZ0\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__8261\,
            I => \N__8256\
        );

    \I__1760\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8252\
        );

    \I__1759\ : InMux
    port map (
            O => \N__8259\,
            I => \N__8246\
        );

    \I__1758\ : InMux
    port map (
            O => \N__8256\,
            I => \N__8243\
        );

    \I__1757\ : InMux
    port map (
            O => \N__8255\,
            I => \N__8240\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__8252\,
            I => \N__8237\
        );

    \I__1755\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8234\
        );

    \I__1754\ : InMux
    port map (
            O => \N__8250\,
            I => \N__8229\
        );

    \I__1753\ : InMux
    port map (
            O => \N__8249\,
            I => \N__8229\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__8246\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__8243\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__8240\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1749\ : Odrv4
    port map (
            O => \N__8237\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1748\ : LocalMux
    port map (
            O => \N__8234\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1747\ : LocalMux
    port map (
            O => \N__8229\,
            I => \U712_REG_SM.C3_SYNCZ0Z_1\
        );

    \I__1746\ : InMux
    port map (
            O => \N__8216\,
            I => \N__8210\
        );

    \I__1745\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8203\
        );

    \I__1744\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8203\
        );

    \I__1743\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8203\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__8210\,
            I => \U712_REG_SM.N_288\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__8203\,
            I => \U712_REG_SM.N_288\
        );

    \I__1740\ : IoInMux
    port map (
            O => \N__8198\,
            I => \N__8195\
        );

    \I__1739\ : LocalMux
    port map (
            O => \N__8195\,
            I => \N__8192\
        );

    \I__1738\ : IoSpan4Mux
    port map (
            O => \N__8192\,
            I => \N__8189\
        );

    \I__1737\ : Sp12to4
    port map (
            O => \N__8189\,
            I => \N__8186\
        );

    \I__1736\ : Span12Mux_s7_v
    port map (
            O => \N__8186\,
            I => \N__8183\
        );

    \I__1735\ : Odrv12
    port map (
            O => \N__8183\,
            I => \CASn_c\
        );

    \I__1734\ : InMux
    port map (
            O => \N__8180\,
            I => \N__8177\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__8177\,
            I => \N__8174\
        );

    \I__1732\ : Odrv4
    port map (
            O => \N__8174\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\
        );

    \I__1731\ : IoInMux
    port map (
            O => \N__8171\,
            I => \N__8168\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__8168\,
            I => \N__8165\
        );

    \I__1729\ : IoSpan4Mux
    port map (
            O => \N__8165\,
            I => \N__8162\
        );

    \I__1728\ : Sp12to4
    port map (
            O => \N__8162\,
            I => \N__8159\
        );

    \I__1727\ : Span12Mux_s3_h
    port map (
            O => \N__8159\,
            I => \N__8156\
        );

    \I__1726\ : Span12Mux_h
    port map (
            O => \N__8156\,
            I => \N__8153\
        );

    \I__1725\ : Odrv12
    port map (
            O => \N__8153\,
            I => \CMA_c_7\
        );

    \I__1724\ : InMux
    port map (
            O => \N__8150\,
            I => \N__8147\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__8147\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\
        );

    \I__1722\ : InMux
    port map (
            O => \N__8144\,
            I => \N__8141\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__8141\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\
        );

    \I__1720\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8135\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__8135\,
            I => \N__8132\
        );

    \I__1718\ : Odrv12
    port map (
            O => \N__8132\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\
        );

    \I__1717\ : InMux
    port map (
            O => \N__8129\,
            I => \N__8126\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8123\
        );

    \I__1715\ : Odrv12
    port map (
            O => \N__8123\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\
        );

    \I__1714\ : InMux
    port map (
            O => \N__8120\,
            I => \N__8117\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__8117\,
            I => \N__8114\
        );

    \I__1712\ : Span4Mux_h
    port map (
            O => \N__8114\,
            I => \N__8111\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__8111\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\
        );

    \I__1710\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8105\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__8105\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__8102\,
            I => \N__8099\
        );

    \I__1707\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8096\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__8096\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\
        );

    \I__1705\ : InMux
    port map (
            O => \N__8093\,
            I => \N__8090\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__8090\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\
        );

    \I__1703\ : InMux
    port map (
            O => \N__8087\,
            I => \N__8080\
        );

    \I__1702\ : InMux
    port map (
            O => \N__8086\,
            I => \N__8077\
        );

    \I__1701\ : InMux
    port map (
            O => \N__8085\,
            I => \N__8073\
        );

    \I__1700\ : InMux
    port map (
            O => \N__8084\,
            I => \N__8068\
        );

    \I__1699\ : InMux
    port map (
            O => \N__8083\,
            I => \N__8068\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__8080\,
            I => \N__8063\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__8077\,
            I => \N__8063\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8076\,
            I => \N__8060\
        );

    \I__1695\ : LocalMux
    port map (
            O => \N__8073\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8068\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__8063\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__8060\,
            I => \U712_REG_SM.LATCH_REG_0_sqmuxa\
        );

    \I__1691\ : IoInMux
    port map (
            O => \N__8051\,
            I => \N__8048\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__8048\,
            I => \N__8045\
        );

    \I__1689\ : Span4Mux_s1_v
    port map (
            O => \N__8045\,
            I => \N__8041\
        );

    \I__1688\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1687\ : Sp12to4
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1685\ : Span12Mux_h
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1684\ : Span4Mux_v
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1683\ : Span12Mux_v
    port map (
            O => \N__8029\,
            I => \N__8021\
        );

    \I__1682\ : Sp12to4
    port map (
            O => \N__8026\,
            I => \N__8021\
        );

    \I__1681\ : Span12Mux_h
    port map (
            O => \N__8021\,
            I => \N__8018\
        );

    \I__1680\ : Span12Mux_v
    port map (
            O => \N__8018\,
            I => \N__8015\
        );

    \I__1679\ : Odrv12
    port map (
            O => \N__8015\,
            I => \RAMENn_c\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8012\,
            I => \N__8008\
        );

    \I__1677\ : InMux
    port map (
            O => \N__8011\,
            I => \N__8005\
        );

    \I__1676\ : InMux
    port map (
            O => \N__8008\,
            I => \N__8002\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__8005\,
            I => \N__7999\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__7999\,
            I => \N__7993\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__7996\,
            I => \N__7990\
        );

    \I__1671\ : Span4Mux_h
    port map (
            O => \N__7993\,
            I => \N__7987\
        );

    \I__1670\ : Sp12to4
    port map (
            O => \N__7990\,
            I => \N__7984\
        );

    \I__1669\ : Sp12to4
    port map (
            O => \N__7987\,
            I => \N__7981\
        );

    \I__1668\ : Span12Mux_h
    port map (
            O => \N__7984\,
            I => \N__7978\
        );

    \I__1667\ : Span12Mux_v
    port map (
            O => \N__7981\,
            I => \N__7975\
        );

    \I__1666\ : Odrv12
    port map (
            O => \N__7978\,
            I => \TSn_c\
        );

    \I__1665\ : Odrv12
    port map (
            O => \N__7975\,
            I => \TSn_c\
        );

    \I__1664\ : InMux
    port map (
            O => \N__7970\,
            I => \N__7964\
        );

    \I__1663\ : InMux
    port map (
            O => \N__7969\,
            I => \N__7964\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7964\,
            I => \U712_REG_SM.CYCLE_RUNZ0\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7961\,
            I => \N__7958\
        );

    \I__1660\ : LocalMux
    port map (
            O => \N__7958\,
            I => \N__7954\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7957\,
            I => \N__7951\
        );

    \I__1658\ : Span4Mux_h
    port map (
            O => \N__7954\,
            I => \N__7947\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__7951\,
            I => \N__7944\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7950\,
            I => \N__7941\
        );

    \I__1655\ : Odrv4
    port map (
            O => \N__7947\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1654\ : Odrv4
    port map (
            O => \N__7944\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7941\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_1\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7931\
        );

    \I__1651\ : LocalMux
    port map (
            O => \N__7931\,
            I => \N__7928\
        );

    \I__1650\ : Span4Mux_v
    port map (
            O => \N__7928\,
            I => \N__7923\
        );

    \I__1649\ : InMux
    port map (
            O => \N__7927\,
            I => \N__7920\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__7926\,
            I => \N__7916\
        );

    \I__1647\ : Span4Mux_v
    port map (
            O => \N__7923\,
            I => \N__7913\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7920\,
            I => \N__7910\
        );

    \I__1645\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7905\
        );

    \I__1644\ : InMux
    port map (
            O => \N__7916\,
            I => \N__7905\
        );

    \I__1643\ : Span4Mux_v
    port map (
            O => \N__7913\,
            I => \N__7900\
        );

    \I__1642\ : Span4Mux_v
    port map (
            O => \N__7910\,
            I => \N__7900\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__7905\,
            I => \N__7897\
        );

    \I__1640\ : Sp12to4
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__1639\ : Span12Mux_v
    port map (
            O => \N__7897\,
            I => \N__7891\
        );

    \I__1638\ : Span12Mux_h
    port map (
            O => \N__7894\,
            I => \N__7888\
        );

    \I__1637\ : Span12Mux_h
    port map (
            O => \N__7891\,
            I => \N__7885\
        );

    \I__1636\ : Odrv12
    port map (
            O => \N__7888\,
            I => \RnW_c\
        );

    \I__1635\ : Odrv12
    port map (
            O => \N__7885\,
            I => \RnW_c\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7880\,
            I => \N__7876\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \N__7870\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__7876\,
            I => \N__7867\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7875\,
            I => \N__7862\
        );

    \I__1630\ : InMux
    port map (
            O => \N__7874\,
            I => \N__7862\
        );

    \I__1629\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7859\
        );

    \I__1628\ : InMux
    port map (
            O => \N__7870\,
            I => \N__7856\
        );

    \I__1627\ : Span4Mux_v
    port map (
            O => \N__7867\,
            I => \N__7851\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__7862\,
            I => \N__7851\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__7859\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__7856\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1623\ : Odrv4
    port map (
            O => \N__7851\,
            I => \REG_WRITE_CYCLE\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__7844\,
            I => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\
        );

    \I__1621\ : IoInMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__7838\,
            I => \N__7835\
        );

    \I__1619\ : Span4Mux_s3_v
    port map (
            O => \N__7835\,
            I => \N__7832\
        );

    \I__1618\ : Span4Mux_v
    port map (
            O => \N__7832\,
            I => \N__7829\
        );

    \I__1617\ : Span4Mux_h
    port map (
            O => \N__7829\,
            I => \N__7826\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__7826\,
            I => \CMA_c_0\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7823\,
            I => \N__7820\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__7820\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\
        );

    \I__1613\ : IoInMux
    port map (
            O => \N__7817\,
            I => \N__7814\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__7814\,
            I => \N__7811\
        );

    \I__1611\ : Span4Mux_s3_v
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1610\ : Span4Mux_v
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1609\ : Span4Mux_v
    port map (
            O => \N__7805\,
            I => \N__7802\
        );

    \I__1608\ : Odrv4
    port map (
            O => \N__7802\,
            I => \CMA_c_2\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7799\,
            I => \N__7795\
        );

    \I__1606\ : InMux
    port map (
            O => \N__7798\,
            I => \N__7792\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__7795\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7792\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\
        );

    \I__1603\ : InMux
    port map (
            O => \N__7787\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\
        );

    \I__1602\ : InMux
    port map (
            O => \N__7784\,
            I => \N__7780\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7777\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__7780\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__7777\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\
        );

    \I__1598\ : InMux
    port map (
            O => \N__7772\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\
        );

    \I__1597\ : InMux
    port map (
            O => \N__7769\,
            I => \N__7765\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7765\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__7762\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__7757\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__7754\,
            I => \N__7750\
        );

    \I__1591\ : InMux
    port map (
            O => \N__7753\,
            I => \N__7747\
        );

    \I__1590\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__7747\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__7744\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\
        );

    \I__1587\ : InMux
    port map (
            O => \N__7739\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\
        );

    \I__1586\ : InMux
    port map (
            O => \N__7736\,
            I => \N__7732\
        );

    \I__1585\ : InMux
    port map (
            O => \N__7735\,
            I => \N__7729\
        );

    \I__1584\ : LocalMux
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7729\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1582\ : Odrv4
    port map (
            O => \N__7726\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\
        );

    \I__1581\ : InMux
    port map (
            O => \N__7721\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7718\,
            I => \N__7714\
        );

    \I__1579\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__1578\ : LocalMux
    port map (
            O => \N__7714\,
            I => \N__7708\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7711\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__7708\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\
        );

    \I__1575\ : InMux
    port map (
            O => \N__7703\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7700\,
            I => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\
        );

    \I__1573\ : InMux
    port map (
            O => \N__7697\,
            I => \N__7694\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7694\,
            I => \N__7690\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7687\
        );

    \I__1570\ : Span4Mux_h
    port map (
            O => \N__7690\,
            I => \N__7684\
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__7687\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1568\ : Odrv4
    port map (
            O => \N__7684\,
            I => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\
        );

    \I__1567\ : ClkMux
    port map (
            O => \N__7679\,
            I => \N__7658\
        );

    \I__1566\ : ClkMux
    port map (
            O => \N__7678\,
            I => \N__7658\
        );

    \I__1565\ : ClkMux
    port map (
            O => \N__7677\,
            I => \N__7658\
        );

    \I__1564\ : ClkMux
    port map (
            O => \N__7676\,
            I => \N__7658\
        );

    \I__1563\ : ClkMux
    port map (
            O => \N__7675\,
            I => \N__7658\
        );

    \I__1562\ : ClkMux
    port map (
            O => \N__7674\,
            I => \N__7658\
        );

    \I__1561\ : ClkMux
    port map (
            O => \N__7673\,
            I => \N__7658\
        );

    \I__1560\ : GlobalMux
    port map (
            O => \N__7658\,
            I => \N__7655\
        );

    \I__1559\ : gio2CtrlBuf
    port map (
            O => \N__7655\,
            I => \C1_c_g\
        );

    \I__1558\ : SRMux
    port map (
            O => \N__7652\,
            I => \N__7649\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7649\,
            I => \N__7646\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__7646\,
            I => \N__7643\
        );

    \I__1555\ : Odrv4
    port map (
            O => \N__7643\,
            I => \U712_CHIP_RAM.REFRESH_RST\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7640\,
            I => \N__7637\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__7637\,
            I => \U712_REG_SM.UDSn_7_iv_i_0_0\
        );

    \I__1552\ : InMux
    port map (
            O => \N__7634\,
            I => \N__7630\
        );

    \I__1551\ : InMux
    port map (
            O => \N__7633\,
            I => \N__7627\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7630\,
            I => \U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__7627\,
            I => \U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1\
        );

    \I__1548\ : InMux
    port map (
            O => \N__7622\,
            I => \N__7619\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__7619\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\
        );

    \I__1546\ : InMux
    port map (
            O => \N__7616\,
            I => \N__7613\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__7613\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\
        );

    \I__1544\ : InMux
    port map (
            O => \N__7610\,
            I => \N__7607\
        );

    \I__1543\ : LocalMux
    port map (
            O => \N__7607\,
            I => \N__7604\
        );

    \I__1542\ : Odrv12
    port map (
            O => \N__7604\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\
        );

    \I__1541\ : InMux
    port map (
            O => \N__7601\,
            I => \N__7598\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__7598\,
            I => \N__7595\
        );

    \I__1539\ : Span12Mux_v
    port map (
            O => \N__7595\,
            I => \N__7592\
        );

    \I__1538\ : Span12Mux_h
    port map (
            O => \N__7592\,
            I => \N__7589\
        );

    \I__1537\ : Odrv12
    port map (
            O => \N__7589\,
            I => \A_c_7\
        );

    \I__1536\ : InMux
    port map (
            O => \N__7586\,
            I => \N__7583\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__7583\,
            I => \U712_CHIP_RAM.N_329\
        );

    \I__1534\ : InMux
    port map (
            O => \N__7580\,
            I => \N__7577\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__7577\,
            I => \N__7574\
        );

    \I__1532\ : Sp12to4
    port map (
            O => \N__7574\,
            I => \N__7571\
        );

    \I__1531\ : Span12Mux_v
    port map (
            O => \N__7571\,
            I => \N__7568\
        );

    \I__1530\ : Span12Mux_h
    port map (
            O => \N__7568\,
            I => \N__7565\
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__7565\,
            I => \A_c_2\
        );

    \I__1528\ : InMux
    port map (
            O => \N__7562\,
            I => \N__7559\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7559\,
            I => \N__7556\
        );

    \I__1526\ : Span12Mux_v
    port map (
            O => \N__7556\,
            I => \N__7553\
        );

    \I__1525\ : Span12Mux_h
    port map (
            O => \N__7553\,
            I => \N__7550\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__7550\,
            I => \A_c_9\
        );

    \I__1523\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7544\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7541\
        );

    \I__1521\ : Span4Mux_h
    port map (
            O => \N__7541\,
            I => \N__7538\
        );

    \I__1520\ : Odrv4
    port map (
            O => \N__7538\,
            I => \U712_CHIP_RAM.REFRESH5lto7_0\
        );

    \I__1519\ : InMux
    port map (
            O => \N__7535\,
            I => \N__7532\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__7532\,
            I => \N__7529\
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__7529\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\
        );

    \I__1516\ : InMux
    port map (
            O => \N__7526\,
            I => \N__7523\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__7523\,
            I => \U712_CHIP_RAM.REFRESH5lto0\
        );

    \I__1514\ : InMux
    port map (
            O => \N__7520\,
            I => \bfn_12_10_0_\
        );

    \I__1513\ : InMux
    port map (
            O => \N__7517\,
            I => \N__7513\
        );

    \I__1512\ : IoInMux
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__7513\,
            I => \N__7507\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7504\
        );

    \I__1509\ : Span4Mux_v
    port map (
            O => \N__7507\,
            I => \N__7501\
        );

    \I__1508\ : IoSpan4Mux
    port map (
            O => \N__7504\,
            I => \N__7498\
        );

    \I__1507\ : Sp12to4
    port map (
            O => \N__7501\,
            I => \N__7495\
        );

    \I__1506\ : IoSpan4Mux
    port map (
            O => \N__7498\,
            I => \N__7492\
        );

    \I__1505\ : Span12Mux_h
    port map (
            O => \N__7495\,
            I => \N__7489\
        );

    \I__1504\ : IoSpan4Mux
    port map (
            O => \N__7492\,
            I => \N__7486\
        );

    \I__1503\ : Odrv12
    port map (
            O => \N__7489\,
            I => \C1_c\
        );

    \I__1502\ : Odrv4
    port map (
            O => \N__7486\,
            I => \C1_c\
        );

    \I__1501\ : InMux
    port map (
            O => \N__7481\,
            I => \N__7478\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__7478\,
            I => \U712_REG_SM.C1_SYNCZ0Z_0\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__7475\,
            I => \N__7472\
        );

    \I__1498\ : InMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1496\ : Odrv4
    port map (
            O => \N__7466\,
            I => \U712_REG_SM.LDSn_7_iv_i_0_0\
        );

    \I__1495\ : InMux
    port map (
            O => \N__7463\,
            I => \N__7460\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__7460\,
            I => \U712_REG_SM.N_278\
        );

    \I__1493\ : IoInMux
    port map (
            O => \N__7457\,
            I => \N__7454\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__7454\,
            I => \N__7451\
        );

    \I__1491\ : IoSpan4Mux
    port map (
            O => \N__7451\,
            I => \N__7448\
        );

    \I__1490\ : Span4Mux_s3_v
    port map (
            O => \N__7448\,
            I => \N__7445\
        );

    \I__1489\ : Sp12to4
    port map (
            O => \N__7445\,
            I => \N__7442\
        );

    \I__1488\ : Span12Mux_s11_v
    port map (
            O => \N__7442\,
            I => \N__7438\
        );

    \I__1487\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__1486\ : Odrv12
    port map (
            O => \N__7438\,
            I => \ASn_c\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__7435\,
            I => \ASn_c\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__7430\,
            I => \N__7427\
        );

    \I__1483\ : InMux
    port map (
            O => \N__7427\,
            I => \N__7423\
        );

    \I__1482\ : InMux
    port map (
            O => \N__7426\,
            I => \N__7420\
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__7423\,
            I => \N__7411\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__7420\,
            I => \N__7411\
        );

    \I__1479\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7407\
        );

    \I__1478\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7401\
        );

    \I__1477\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7401\
        );

    \I__1476\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7398\
        );

    \I__1475\ : Span12Mux_v
    port map (
            O => \N__7411\,
            I => \N__7395\
        );

    \I__1474\ : InMux
    port map (
            O => \N__7410\,
            I => \N__7392\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__7407\,
            I => \N__7389\
        );

    \I__1472\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7386\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__7401\,
            I => \N__7381\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__7398\,
            I => \N__7381\
        );

    \I__1469\ : Odrv12
    port map (
            O => \N__7395\,
            I => \WRITE_CYCLE\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__7392\,
            I => \WRITE_CYCLE\
        );

    \I__1467\ : Odrv4
    port map (
            O => \N__7389\,
            I => \WRITE_CYCLE\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__7386\,
            I => \WRITE_CYCLE\
        );

    \I__1465\ : Odrv4
    port map (
            O => \N__7381\,
            I => \WRITE_CYCLE\
        );

    \I__1464\ : IoInMux
    port map (
            O => \N__7370\,
            I => \N__7367\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__7367\,
            I => \N__7364\
        );

    \I__1462\ : Span4Mux_s0_v
    port map (
            O => \N__7364\,
            I => \N__7361\
        );

    \I__1461\ : Sp12to4
    port map (
            O => \N__7361\,
            I => \N__7358\
        );

    \I__1460\ : Span12Mux_h
    port map (
            O => \N__7358\,
            I => \N__7355\
        );

    \I__1459\ : Odrv12
    port map (
            O => \N__7355\,
            I => \N_259\
        );

    \I__1458\ : IoInMux
    port map (
            O => \N__7352\,
            I => \N__7349\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__7349\,
            I => \N__7346\
        );

    \I__1456\ : IoSpan4Mux
    port map (
            O => \N__7346\,
            I => \N__7343\
        );

    \I__1455\ : Sp12to4
    port map (
            O => \N__7343\,
            I => \N__7340\
        );

    \I__1454\ : Span12Mux_v
    port map (
            O => \N__7340\,
            I => \N__7337\
        );

    \I__1453\ : Span12Mux_h
    port map (
            O => \N__7337\,
            I => \N__7331\
        );

    \I__1452\ : InMux
    port map (
            O => \N__7336\,
            I => \N__7328\
        );

    \I__1451\ : InMux
    port map (
            O => \N__7335\,
            I => \N__7325\
        );

    \I__1450\ : InMux
    port map (
            O => \N__7334\,
            I => \N__7322\
        );

    \I__1449\ : Odrv12
    port map (
            O => \N__7331\,
            I => \LDSn_c\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__7328\,
            I => \LDSn_c\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__7325\,
            I => \LDSn_c\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__7322\,
            I => \LDSn_c\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__7313\,
            I => \U712_REG_SM.N_467_cascade_\
        );

    \I__1444\ : InMux
    port map (
            O => \N__7310\,
            I => \N__7307\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__7307\,
            I => \U712_REG_SM.N_371\
        );

    \I__1442\ : InMux
    port map (
            O => \N__7304\,
            I => \N__7301\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7301\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\
        );

    \I__1440\ : IoInMux
    port map (
            O => \N__7298\,
            I => \N__7295\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__7295\,
            I => \N__7292\
        );

    \I__1438\ : Odrv12
    port map (
            O => \N__7292\,
            I => \CMA_c_1\
        );

    \I__1437\ : InMux
    port map (
            O => \N__7289\,
            I => \N__7286\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7286\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\
        );

    \I__1435\ : InMux
    port map (
            O => \N__7283\,
            I => \N__7280\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__7280\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\
        );

    \I__1433\ : IoInMux
    port map (
            O => \N__7277\,
            I => \N__7274\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__7274\,
            I => \N__7271\
        );

    \I__1431\ : IoSpan4Mux
    port map (
            O => \N__7271\,
            I => \N__7268\
        );

    \I__1430\ : Span4Mux_s2_h
    port map (
            O => \N__7268\,
            I => \N__7265\
        );

    \I__1429\ : Sp12to4
    port map (
            O => \N__7265\,
            I => \N__7262\
        );

    \I__1428\ : Span12Mux_h
    port map (
            O => \N__7262\,
            I => \N__7259\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__7259\,
            I => \CMA_c_5\
        );

    \I__1426\ : InMux
    port map (
            O => \N__7256\,
            I => \N__7253\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__7253\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__7250\,
            I => \N__7247\
        );

    \I__1423\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7244\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__7244\,
            I => \U712_BYTE_ENABLE.N_92\
        );

    \I__1421\ : IoInMux
    port map (
            O => \N__7241\,
            I => \N__7238\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__7238\,
            I => \N__7235\
        );

    \I__1419\ : IoSpan4Mux
    port map (
            O => \N__7235\,
            I => \N__7232\
        );

    \I__1418\ : Span4Mux_s2_h
    port map (
            O => \N__7232\,
            I => \N__7229\
        );

    \I__1417\ : Sp12to4
    port map (
            O => \N__7229\,
            I => \N__7226\
        );

    \I__1416\ : Span12Mux_s9_h
    port map (
            O => \N__7226\,
            I => \N__7223\
        );

    \I__1415\ : Span12Mux_v
    port map (
            O => \N__7223\,
            I => \N__7220\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__7220\,
            I => \N_315\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7217\,
            I => \U712_REG_SM.N_278_cascade_\
        );

    \I__1412\ : CascadeMux
    port map (
            O => \N__7214\,
            I => \N__7210\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__7213\,
            I => \N__7207\
        );

    \I__1410\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7200\
        );

    \I__1409\ : InMux
    port map (
            O => \N__7207\,
            I => \N__7197\
        );

    \I__1408\ : InMux
    port map (
            O => \N__7206\,
            I => \N__7192\
        );

    \I__1407\ : InMux
    port map (
            O => \N__7205\,
            I => \N__7192\
        );

    \I__1406\ : InMux
    port map (
            O => \N__7204\,
            I => \N__7187\
        );

    \I__1405\ : InMux
    port map (
            O => \N__7203\,
            I => \N__7187\
        );

    \I__1404\ : LocalMux
    port map (
            O => \N__7200\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__7197\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__7192\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__7187\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_7\
        );

    \I__1400\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7175\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__7175\,
            I => \N__7171\
        );

    \I__1398\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7168\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__7171\,
            I => \U712_REG_SM.N_272\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__7168\,
            I => \U712_REG_SM.N_272\
        );

    \I__1395\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7157\
        );

    \I__1394\ : InMux
    port map (
            O => \N__7162\,
            I => \N__7157\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__7157\,
            I => \U712_REG_SM.N_309\
        );

    \I__1392\ : CascadeMux
    port map (
            O => \N__7154\,
            I => \U712_REG_SM.N_272_cascade_\
        );

    \I__1391\ : IoInMux
    port map (
            O => \N__7151\,
            I => \N__7148\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__7148\,
            I => \N__7145\
        );

    \I__1389\ : IoSpan4Mux
    port map (
            O => \N__7145\,
            I => \N__7142\
        );

    \I__1388\ : Span4Mux_s3_h
    port map (
            O => \N__7142\,
            I => \N__7139\
        );

    \I__1387\ : Span4Mux_h
    port map (
            O => \N__7139\,
            I => \N__7136\
        );

    \I__1386\ : Sp12to4
    port map (
            O => \N__7136\,
            I => \N__7133\
        );

    \I__1385\ : Span12Mux_h
    port map (
            O => \N__7133\,
            I => \N__7129\
        );

    \I__1384\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7126\
        );

    \I__1383\ : Span12Mux_h
    port map (
            O => \N__7129\,
            I => \N__7123\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__7126\,
            I => \N__7120\
        );

    \I__1381\ : Span12Mux_v
    port map (
            O => \N__7123\,
            I => \N__7117\
        );

    \I__1380\ : Span12Mux_h
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1379\ : Odrv12
    port map (
            O => \N__7117\,
            I => \C3_c\
        );

    \I__1378\ : Odrv12
    port map (
            O => \N__7114\,
            I => \C3_c\
        );

    \I__1377\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7106\
        );

    \I__1376\ : LocalMux
    port map (
            O => \N__7106\,
            I => \U712_REG_SM.C3_SYNCZ0Z_0\
        );

    \I__1375\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7100\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__7100\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\
        );

    \I__1373\ : InMux
    port map (
            O => \N__7097\,
            I => \N__7091\
        );

    \I__1372\ : InMux
    port map (
            O => \N__7096\,
            I => \N__7091\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__7091\,
            I => \N__7088\
        );

    \I__1370\ : Span4Mux_v
    port map (
            O => \N__7088\,
            I => \N__7085\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__7085\,
            I => \N__7082\
        );

    \I__1368\ : Sp12to4
    port map (
            O => \N__7082\,
            I => \N__7079\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__7079\,
            I => \N__7076\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__7076\,
            I => \A_c_14\
        );

    \I__1365\ : InMux
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__7070\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\
        );

    \I__1363\ : InMux
    port map (
            O => \N__7067\,
            I => \N__7064\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7064\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\
        );

    \I__1361\ : InMux
    port map (
            O => \N__7061\,
            I => \N__7058\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__7058\,
            I => \N__7055\
        );

    \I__1359\ : Odrv4
    port map (
            O => \N__7055\,
            I => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\
        );

    \I__1358\ : IoInMux
    port map (
            O => \N__7052\,
            I => \N__7049\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__7049\,
            I => \N__7046\
        );

    \I__1356\ : Span4Mux_s2_v
    port map (
            O => \N__7046\,
            I => \N__7043\
        );

    \I__1355\ : Span4Mux_h
    port map (
            O => \N__7043\,
            I => \N__7040\
        );

    \I__1354\ : Sp12to4
    port map (
            O => \N__7040\,
            I => \N__7036\
        );

    \I__1353\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7033\
        );

    \I__1352\ : Span12Mux_v
    port map (
            O => \N__7036\,
            I => \N__7026\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__7033\,
            I => \N__7026\
        );

    \I__1350\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7023\
        );

    \I__1349\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7020\
        );

    \I__1348\ : Odrv12
    port map (
            O => \N__7026\,
            I => \DBENn_c\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__7023\,
            I => \DBENn_c\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__7020\,
            I => \DBENn_c\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7013\,
            I => \N__7009\
        );

    \I__1344\ : InMux
    port map (
            O => \N__7012\,
            I => \N__7005\
        );

    \I__1343\ : InMux
    port map (
            O => \N__7009\,
            I => \N__7002\
        );

    \I__1342\ : InMux
    port map (
            O => \N__7008\,
            I => \N__6997\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__7005\,
            I => \N__6994\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__7002\,
            I => \N__6991\
        );

    \I__1339\ : InMux
    port map (
            O => \N__7001\,
            I => \N__6988\
        );

    \I__1338\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6984\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__6997\,
            I => \N__6981\
        );

    \I__1336\ : Span4Mux_v
    port map (
            O => \N__6994\,
            I => \N__6976\
        );

    \I__1335\ : Span4Mux_v
    port map (
            O => \N__6991\,
            I => \N__6976\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6988\,
            I => \N__6973\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6970\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6984\,
            I => \N__6967\
        );

    \I__1331\ : Odrv12
    port map (
            O => \N__6981\,
            I => \DMA_CYCLE\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__6976\,
            I => \DMA_CYCLE\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__6973\,
            I => \DMA_CYCLE\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__6970\,
            I => \DMA_CYCLE\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__6967\,
            I => \DMA_CYCLE\
        );

    \I__1326\ : InMux
    port map (
            O => \N__6956\,
            I => \N__6953\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6953\,
            I => \N__6950\
        );

    \I__1324\ : Span4Mux_h
    port map (
            O => \N__6950\,
            I => \N__6947\
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6947\,
            I => \U712_CHIP_RAM.REFRESH5lt7\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6940\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6940\,
            I => \N__6932\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6932\
        );

    \I__1318\ : Odrv12
    port map (
            O => \N__6932\,
            I => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\
        );

    \I__1317\ : IoInMux
    port map (
            O => \N__6929\,
            I => \N__6926\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6926\,
            I => \N__6923\
        );

    \I__1315\ : IoSpan4Mux
    port map (
            O => \N__6923\,
            I => \N__6920\
        );

    \I__1314\ : Span4Mux_s3_h
    port map (
            O => \N__6920\,
            I => \N__6917\
        );

    \I__1313\ : Sp12to4
    port map (
            O => \N__6917\,
            I => \N__6914\
        );

    \I__1312\ : Span12Mux_h
    port map (
            O => \N__6914\,
            I => \N__6911\
        );

    \I__1311\ : Span12Mux_v
    port map (
            O => \N__6911\,
            I => \N__6908\
        );

    \I__1310\ : Odrv12
    port map (
            O => \N__6908\,
            I => \N_49_i\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6905\,
            I => \N__6899\
        );

    \I__1308\ : InMux
    port map (
            O => \N__6904\,
            I => \N__6899\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__6899\,
            I => \U712_REG_SM.STATE_COUNTERc_0\
        );

    \I__1306\ : InMux
    port map (
            O => \N__6896\,
            I => \N__6893\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6893\,
            I => \U712_REG_SM.un15_0_i_0_0\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__6890\,
            I => \N__6887\
        );

    \I__1303\ : InMux
    port map (
            O => \N__6887\,
            I => \N__6884\
        );

    \I__1302\ : LocalMux
    port map (
            O => \N__6884\,
            I => \U712_REG_SM.N_297\
        );

    \I__1301\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6875\
        );

    \I__1300\ : InMux
    port map (
            O => \N__6880\,
            I => \N__6872\
        );

    \I__1299\ : InMux
    port map (
            O => \N__6879\,
            I => \N__6869\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6866\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6875\,
            I => \N__6862\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__6872\,
            I => \N__6857\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__6869\,
            I => \N__6857\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6854\
        );

    \I__1293\ : InMux
    port map (
            O => \N__6865\,
            I => \N__6851\
        );

    \I__1292\ : Span4Mux_v
    port map (
            O => \N__6862\,
            I => \N__6848\
        );

    \I__1291\ : Span4Mux_h
    port map (
            O => \N__6857\,
            I => \N__6843\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__6854\,
            I => \N__6843\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6851\,
            I => \REG_TACK\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__6848\,
            I => \REG_TACK\
        );

    \I__1287\ : Odrv4
    port map (
            O => \N__6843\,
            I => \REG_TACK\
        );

    \I__1286\ : InMux
    port map (
            O => \N__6836\,
            I => \N__6831\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6835\,
            I => \N__6828\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6834\,
            I => \N__6825\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6831\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6828\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6825\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_6\
        );

    \I__1280\ : IoInMux
    port map (
            O => \N__6818\,
            I => \N__6815\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__6815\,
            I => \N__6812\
        );

    \I__1278\ : Span12Mux_s11_v
    port map (
            O => \N__6812\,
            I => \N__6808\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6811\,
            I => \N__6805\
        );

    \I__1276\ : Odrv12
    port map (
            O => \N__6808\,
            I => \REGENn_c\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6805\,
            I => \REGENn_c\
        );

    \I__1274\ : InMux
    port map (
            O => \N__6800\,
            I => \N__6793\
        );

    \I__1273\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6793\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6790\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6793\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__6790\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_4\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__6785\,
            I => \N__6781\
        );

    \I__1268\ : InMux
    port map (
            O => \N__6784\,
            I => \N__6777\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6781\,
            I => \N__6774\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6780\,
            I => \N__6771\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6777\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6774\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__6771\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_3\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6764\,
            I => \N__6761\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__6761\,
            I => \N__6757\
        );

    \I__1260\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6754\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__6757\,
            I => \N__6748\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__6754\,
            I => \N__6748\
        );

    \I__1257\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6745\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__6748\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6745\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_1\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__6740\,
            I => \N__6731\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6739\,
            I => \N__6726\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6738\,
            I => \N__6721\
        );

    \I__1251\ : InMux
    port map (
            O => \N__6737\,
            I => \N__6721\
        );

    \I__1250\ : InMux
    port map (
            O => \N__6736\,
            I => \N__6716\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6735\,
            I => \N__6711\
        );

    \I__1248\ : InMux
    port map (
            O => \N__6734\,
            I => \N__6711\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6731\,
            I => \N__6708\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6730\,
            I => \N__6703\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6729\,
            I => \N__6703\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__6726\,
            I => \N__6698\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6721\,
            I => \N__6698\
        );

    \I__1242\ : InMux
    port map (
            O => \N__6720\,
            I => \N__6695\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__6719\,
            I => \N__6689\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6716\,
            I => \N__6682\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__6711\,
            I => \N__6682\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6708\,
            I => \N__6677\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__6703\,
            I => \N__6677\
        );

    \I__1236\ : Span4Mux_h
    port map (
            O => \N__6698\,
            I => \N__6672\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6695\,
            I => \N__6672\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6694\,
            I => \N__6665\
        );

    \I__1233\ : InMux
    port map (
            O => \N__6693\,
            I => \N__6665\
        );

    \I__1232\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6665\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6689\,
            I => \N__6660\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6688\,
            I => \N__6660\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6687\,
            I => \N__6657\
        );

    \I__1228\ : Odrv4
    port map (
            O => \N__6682\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1227\ : Odrv12
    port map (
            O => \N__6677\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1226\ : Odrv4
    port map (
            O => \N__6672\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6665\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__6660\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6657\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__6644\,
            I => \U712_CHIP_RAM.N_316_cascade_\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6638\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__6632\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1\
        );

    \I__1217\ : CascadeMux
    port map (
            O => \N__6629\,
            I => \N__6623\
        );

    \I__1216\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6614\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__6627\,
            I => \N__6610\
        );

    \I__1214\ : InMux
    port map (
            O => \N__6626\,
            I => \N__6607\
        );

    \I__1213\ : InMux
    port map (
            O => \N__6623\,
            I => \N__6603\
        );

    \I__1212\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6600\
        );

    \I__1211\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6592\
        );

    \I__1210\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6592\
        );

    \I__1209\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6592\
        );

    \I__1208\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6589\
        );

    \I__1207\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6586\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__6614\,
            I => \N__6583\
        );

    \I__1205\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6578\
        );

    \I__1204\ : InMux
    port map (
            O => \N__6610\,
            I => \N__6575\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6572\
        );

    \I__1202\ : CascadeMux
    port map (
            O => \N__6606\,
            I => \N__6568\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__6603\,
            I => \N__6562\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6562\
        );

    \I__1199\ : InMux
    port map (
            O => \N__6599\,
            I => \N__6559\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N__6554\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6554\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6551\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__6583\,
            I => \N__6548\
        );

    \I__1194\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6543\
        );

    \I__1193\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6543\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__6578\,
            I => \N__6536\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__6575\,
            I => \N__6536\
        );

    \I__1190\ : Span4Mux_h
    port map (
            O => \N__6572\,
            I => \N__6536\
        );

    \I__1189\ : InMux
    port map (
            O => \N__6571\,
            I => \N__6533\
        );

    \I__1188\ : InMux
    port map (
            O => \N__6568\,
            I => \N__6530\
        );

    \I__1187\ : InMux
    port map (
            O => \N__6567\,
            I => \N__6527\
        );

    \I__1186\ : Span4Mux_v
    port map (
            O => \N__6562\,
            I => \N__6518\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__6559\,
            I => \N__6518\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__6554\,
            I => \N__6518\
        );

    \I__1183\ : Span4Mux_h
    port map (
            O => \N__6551\,
            I => \N__6518\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__6548\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__6543\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__6536\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__6533\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__6530\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__6527\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__6518\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\
        );

    \I__1175\ : InMux
    port map (
            O => \N__6503\,
            I => \N__6500\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__6500\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__6497\,
            I => \N__6491\
        );

    \I__1172\ : InMux
    port map (
            O => \N__6496\,
            I => \N__6482\
        );

    \I__1171\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6482\
        );

    \I__1170\ : InMux
    port map (
            O => \N__6494\,
            I => \N__6482\
        );

    \I__1169\ : InMux
    port map (
            O => \N__6491\,
            I => \N__6479\
        );

    \I__1168\ : InMux
    port map (
            O => \N__6490\,
            I => \N__6476\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6489\,
            I => \N__6468\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__6482\,
            I => \N__6461\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6461\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__6476\,
            I => \N__6461\
        );

    \I__1163\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6456\
        );

    \I__1162\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6456\
        );

    \I__1161\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6453\
        );

    \I__1160\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6450\
        );

    \I__1159\ : InMux
    port map (
            O => \N__6471\,
            I => \N__6447\
        );

    \I__1158\ : InMux
    port map (
            O => \N__6468\,
            I => \N__6442\
        );

    \I__1157\ : Span4Mux_v
    port map (
            O => \N__6461\,
            I => \N__6439\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__6456\,
            I => \N__6430\
        );

    \I__1155\ : LocalMux
    port map (
            O => \N__6453\,
            I => \N__6430\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__6450\,
            I => \N__6430\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__6447\,
            I => \N__6430\
        );

    \I__1152\ : InMux
    port map (
            O => \N__6446\,
            I => \N__6425\
        );

    \I__1151\ : InMux
    port map (
            O => \N__6445\,
            I => \N__6425\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__6442\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1149\ : Odrv4
    port map (
            O => \N__6439\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1148\ : Odrv4
    port map (
            O => \N__6430\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6425\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\
        );

    \I__1146\ : CascadeMux
    port map (
            O => \N__6416\,
            I => \N__6412\
        );

    \I__1145\ : CascadeMux
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1144\ : InMux
    port map (
            O => \N__6412\,
            I => \N__6398\
        );

    \I__1143\ : InMux
    port map (
            O => \N__6409\,
            I => \N__6398\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6408\,
            I => \N__6393\
        );

    \I__1141\ : InMux
    port map (
            O => \N__6407\,
            I => \N__6393\
        );

    \I__1140\ : CascadeMux
    port map (
            O => \N__6406\,
            I => \N__6390\
        );

    \I__1139\ : CascadeMux
    port map (
            O => \N__6405\,
            I => \N__6385\
        );

    \I__1138\ : CascadeMux
    port map (
            O => \N__6404\,
            I => \N__6382\
        );

    \I__1137\ : InMux
    port map (
            O => \N__6403\,
            I => \N__6379\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6374\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__6393\,
            I => \N__6374\
        );

    \I__1134\ : InMux
    port map (
            O => \N__6390\,
            I => \N__6367\
        );

    \I__1133\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6364\
        );

    \I__1132\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6361\
        );

    \I__1131\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6355\
        );

    \I__1130\ : InMux
    port map (
            O => \N__6382\,
            I => \N__6352\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6349\
        );

    \I__1128\ : Span4Mux_v
    port map (
            O => \N__6374\,
            I => \N__6346\
        );

    \I__1127\ : InMux
    port map (
            O => \N__6373\,
            I => \N__6341\
        );

    \I__1126\ : InMux
    port map (
            O => \N__6372\,
            I => \N__6341\
        );

    \I__1125\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6336\
        );

    \I__1124\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6336\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__6367\,
            I => \N__6329\
        );

    \I__1122\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6329\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__6361\,
            I => \N__6329\
        );

    \I__1120\ : InMux
    port map (
            O => \N__6360\,
            I => \N__6322\
        );

    \I__1119\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6322\
        );

    \I__1118\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6322\
        );

    \I__1117\ : LocalMux
    port map (
            O => \N__6355\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__6352\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1115\ : Odrv4
    port map (
            O => \N__6349\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1114\ : Odrv4
    port map (
            O => \N__6346\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__6341\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__6336\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1111\ : Odrv4
    port map (
            O => \N__6329\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__6322\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\
        );

    \I__1109\ : InMux
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__6302\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\
        );

    \I__1107\ : InMux
    port map (
            O => \N__6299\,
            I => \N__6290\
        );

    \I__1106\ : InMux
    port map (
            O => \N__6298\,
            I => \N__6287\
        );

    \I__1105\ : InMux
    port map (
            O => \N__6297\,
            I => \N__6282\
        );

    \I__1104\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6282\
        );

    \I__1103\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6277\
        );

    \I__1102\ : InMux
    port map (
            O => \N__6294\,
            I => \N__6277\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__6293\,
            I => \N__6273\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6270\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__6287\,
            I => \N__6259\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__6282\,
            I => \N__6259\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__6277\,
            I => \N__6259\
        );

    \I__1096\ : InMux
    port map (
            O => \N__6276\,
            I => \N__6256\
        );

    \I__1095\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6253\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__6270\,
            I => \N__6250\
        );

    \I__1093\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6245\
        );

    \I__1092\ : InMux
    port map (
            O => \N__6268\,
            I => \N__6245\
        );

    \I__1091\ : InMux
    port map (
            O => \N__6267\,
            I => \N__6240\
        );

    \I__1090\ : InMux
    port map (
            O => \N__6266\,
            I => \N__6240\
        );

    \I__1089\ : Sp12to4
    port map (
            O => \N__6259\,
            I => \N__6235\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6235\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__6253\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1086\ : Odrv4
    port map (
            O => \N__6250\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__6245\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__6240\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1083\ : Odrv12
    port map (
            O => \N__6235\,
            I => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\
        );

    \I__1082\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6218\
        );

    \I__1081\ : InMux
    port map (
            O => \N__6223\,
            I => \N__6215\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__6222\,
            I => \N__6208\
        );

    \I__1079\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6204\
        );

    \I__1078\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6197\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__6215\,
            I => \N__6189\
        );

    \I__1076\ : InMux
    port map (
            O => \N__6214\,
            I => \N__6184\
        );

    \I__1075\ : InMux
    port map (
            O => \N__6213\,
            I => \N__6184\
        );

    \I__1074\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6181\
        );

    \I__1073\ : InMux
    port map (
            O => \N__6211\,
            I => \N__6176\
        );

    \I__1072\ : InMux
    port map (
            O => \N__6208\,
            I => \N__6176\
        );

    \I__1071\ : InMux
    port map (
            O => \N__6207\,
            I => \N__6173\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__6204\,
            I => \N__6170\
        );

    \I__1069\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6165\
        );

    \I__1068\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6165\
        );

    \I__1067\ : InMux
    port map (
            O => \N__6201\,
            I => \N__6162\
        );

    \I__1066\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6157\
        );

    \I__1065\ : Span4Mux_v
    port map (
            O => \N__6197\,
            I => \N__6154\
        );

    \I__1064\ : InMux
    port map (
            O => \N__6196\,
            I => \N__6147\
        );

    \I__1063\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6147\
        );

    \I__1062\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6147\
        );

    \I__1061\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6142\
        );

    \I__1060\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6142\
        );

    \I__1059\ : Span4Mux_v
    port map (
            O => \N__6189\,
            I => \N__6133\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__6184\,
            I => \N__6133\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__6181\,
            I => \N__6133\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__6176\,
            I => \N__6133\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__6173\,
            I => \N__6124\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__6170\,
            I => \N__6124\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__6165\,
            I => \N__6124\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6124\
        );

    \I__1051\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6121\
        );

    \I__1050\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6118\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__6157\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1048\ : Odrv4
    port map (
            O => \N__6154\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__6147\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__6142\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__6133\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__6124\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__6121\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__6118\,
            I => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\
        );

    \I__1041\ : CascadeMux
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1040\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6090\
        );

    \I__1039\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6087\
        );

    \I__1038\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6084\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__6095\,
            I => \N__6081\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__6094\,
            I => \N__6078\
        );

    \I__1035\ : InMux
    port map (
            O => \N__6093\,
            I => \N__6073\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__6090\,
            I => \N__6070\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__6087\,
            I => \N__6067\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__6084\,
            I => \N__6064\
        );

    \I__1031\ : InMux
    port map (
            O => \N__6081\,
            I => \N__6057\
        );

    \I__1030\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6057\
        );

    \I__1029\ : InMux
    port map (
            O => \N__6077\,
            I => \N__6057\
        );

    \I__1028\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6054\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__6073\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1026\ : Odrv4
    port map (
            O => \N__6070\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__6067\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1024\ : Odrv4
    port map (
            O => \N__6064\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__6057\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__6054\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15\
        );

    \I__1021\ : InMux
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__6038\,
            I => \U712_CHIP_RAM.N_109_i\
        );

    \I__1019\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6032\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__6032\,
            I => \N__6029\
        );

    \I__1017\ : Span12Mux_s11_v
    port map (
            O => \N__6029\,
            I => \N__6026\
        );

    \I__1016\ : Span12Mux_h
    port map (
            O => \N__6026\,
            I => \N__6023\
        );

    \I__1015\ : Odrv12
    port map (
            O => \N__6023\,
            I => \A_c_10\
        );

    \I__1014\ : InMux
    port map (
            O => \N__6020\,
            I => \N__6017\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__6017\,
            I => \N__6014\
        );

    \I__1012\ : Span12Mux_v
    port map (
            O => \N__6014\,
            I => \N__6011\
        );

    \I__1011\ : Span12Mux_h
    port map (
            O => \N__6011\,
            I => \N__6008\
        );

    \I__1010\ : Odrv12
    port map (
            O => \N__6008\,
            I => \A_c_16\
        );

    \I__1009\ : InMux
    port map (
            O => \N__6005\,
            I => \N__6002\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__6002\,
            I => \N__5999\
        );

    \I__1007\ : Span12Mux_v
    port map (
            O => \N__5999\,
            I => \N__5996\
        );

    \I__1006\ : Span12Mux_h
    port map (
            O => \N__5996\,
            I => \N__5993\
        );

    \I__1005\ : Odrv12
    port map (
            O => \N__5993\,
            I => \A_c_18\
        );

    \I__1004\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5987\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5987\,
            I => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\
        );

    \I__1002\ : CascadeMux
    port map (
            O => \N__5984\,
            I => \U712_CHIP_RAM.N_411_cascade_\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5981\,
            I => \N__5978\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5978\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__5975\,
            I => \N__5971\
        );

    \I__998\ : CascadeMux
    port map (
            O => \N__5974\,
            I => \N__5967\
        );

    \I__997\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5960\
        );

    \I__996\ : InMux
    port map (
            O => \N__5970\,
            I => \N__5960\
        );

    \I__995\ : InMux
    port map (
            O => \N__5967\,
            I => \N__5960\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5960\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__5957\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_\
        );

    \I__992\ : InMux
    port map (
            O => \N__5954\,
            I => \N__5948\
        );

    \I__991\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5941\
        );

    \I__990\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5941\
        );

    \I__989\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5941\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5948\,
            I => \U712_CHIP_RAM.N_294\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5941\,
            I => \U712_CHIP_RAM.N_294\
        );

    \I__986\ : CEMux
    port map (
            O => \N__5936\,
            I => \N__5932\
        );

    \I__985\ : CEMux
    port map (
            O => \N__5935\,
            I => \N__5929\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5932\,
            I => \N__5926\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__982\ : Span4Mux_v
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__981\ : Span4Mux_h
    port map (
            O => \N__5923\,
            I => \N__5917\
        );

    \I__980\ : Odrv4
    port map (
            O => \N__5920\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__979\ : Odrv4
    port map (
            O => \N__5917\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\
        );

    \I__978\ : InMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__5909\,
            I => \N__5901\
        );

    \I__976\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5897\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__5907\,
            I => \N__5894\
        );

    \I__974\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5888\
        );

    \I__973\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5885\
        );

    \I__972\ : InMux
    port map (
            O => \N__5904\,
            I => \N__5882\
        );

    \I__971\ : Span4Mux_h
    port map (
            O => \N__5901\,
            I => \N__5879\
        );

    \I__970\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5876\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5897\,
            I => \N__5873\
        );

    \I__968\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5870\
        );

    \I__967\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5863\
        );

    \I__966\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5863\
        );

    \I__965\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5863\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5888\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__5885\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5882\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__961\ : Odrv4
    port map (
            O => \N__5879\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5876\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__959\ : Odrv4
    port map (
            O => \N__5873\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5870\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__5863\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\
        );

    \I__956\ : InMux
    port map (
            O => \N__5846\,
            I => \N__5843\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5843\,
            I => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\
        );

    \I__954\ : CascadeMux
    port map (
            O => \N__5840\,
            I => \N__5836\
        );

    \I__953\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \N__5829\
        );

    \I__952\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5826\
        );

    \I__951\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5823\
        );

    \I__950\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5818\
        );

    \I__949\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5818\
        );

    \I__948\ : InMux
    port map (
            O => \N__5832\,
            I => \N__5813\
        );

    \I__947\ : InMux
    port map (
            O => \N__5829\,
            I => \N__5813\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__5826\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__5823\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5818\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5813\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\
        );

    \I__942\ : CascadeMux
    port map (
            O => \N__5804\,
            I => \N__5801\
        );

    \I__941\ : InMux
    port map (
            O => \N__5801\,
            I => \N__5797\
        );

    \I__940\ : InMux
    port map (
            O => \N__5800\,
            I => \N__5794\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5797\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__5794\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\
        );

    \I__937\ : InMux
    port map (
            O => \N__5789\,
            I => \N__5785\
        );

    \I__936\ : InMux
    port map (
            O => \N__5788\,
            I => \N__5781\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__5785\,
            I => \N__5778\
        );

    \I__934\ : InMux
    port map (
            O => \N__5784\,
            I => \N__5775\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5781\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__932\ : Odrv4
    port map (
            O => \N__5778\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5775\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\
        );

    \I__930\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__5765\,
            I => \U712_REG_SM.STATE_COUNTERZ0Z_5\
        );

    \I__928\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5759\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__5759\,
            I => \N__5756\
        );

    \I__926\ : Span4Mux_v
    port map (
            O => \N__5756\,
            I => \N__5752\
        );

    \I__925\ : InMux
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__5752\,
            I => \LATCH_REG\
        );

    \I__923\ : LocalMux
    port map (
            O => \N__5749\,
            I => \LATCH_REG\
        );

    \I__922\ : InMux
    port map (
            O => \N__5744\,
            I => \N__5741\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__5741\,
            I => \N__5738\
        );

    \I__920\ : Span12Mux_v
    port map (
            O => \N__5738\,
            I => \N__5734\
        );

    \I__919\ : InMux
    port map (
            O => \N__5737\,
            I => \N__5731\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__5734\,
            I => \REG_CPU_CYCLE\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5731\,
            I => \REG_CPU_CYCLE\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5726\,
            I => \U712_REG_SM.STATE_COUNTERc_0_cascade_\
        );

    \I__915\ : InMux
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__5720\,
            I => \U712_REG_SM.REG_CPU_CYCLE_e_1\
        );

    \I__913\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5714\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5711\
        );

    \I__911\ : Span12Mux_v
    port map (
            O => \N__5711\,
            I => \N__5708\
        );

    \I__910\ : Span12Mux_h
    port map (
            O => \N__5708\,
            I => \N__5705\
        );

    \I__909\ : Span12Mux_v
    port map (
            O => \N__5705\,
            I => \N__5702\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5702\,
            I => \A_c_3\
        );

    \I__907\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5693\
        );

    \I__906\ : InMux
    port map (
            O => \N__5698\,
            I => \N__5693\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__904\ : Odrv4
    port map (
            O => \N__5690\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__5687\,
            I => \U712_CHIP_RAM.N_421_cascade_\
        );

    \I__902\ : CEMux
    port map (
            O => \N__5684\,
            I => \N__5681\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5681\,
            I => \N__5677\
        );

    \I__900\ : CEMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__899\ : Span4Mux_h
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__897\ : Odrv4
    port map (
            O => \N__5671\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__896\ : Odrv12
    port map (
            O => \N__5668\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\
        );

    \I__895\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5659\
        );

    \I__894\ : InMux
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5659\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5656\,
            I => \U712_CHIP_RAM.DMA_AZ0Z20\
        );

    \I__891\ : InMux
    port map (
            O => \N__5651\,
            I => \N__5648\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5648\,
            I => \U712_CHIP_RAM.N_18\
        );

    \I__889\ : CEMux
    port map (
            O => \N__5645\,
            I => \N__5642\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5642\,
            I => \U712_CHIP_RAM.N_18_0\
        );

    \I__887\ : InMux
    port map (
            O => \N__5639\,
            I => \N__5635\
        );

    \I__886\ : InMux
    port map (
            O => \N__5638\,
            I => \N__5632\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__5632\,
            I => \N__5626\
        );

    \I__883\ : Span4Mux_h
    port map (
            O => \N__5629\,
            I => \N__5623\
        );

    \I__882\ : Odrv4
    port map (
            O => \N__5626\,
            I => \U712_CHIP_RAM.N_113\
        );

    \I__881\ : Odrv4
    port map (
            O => \N__5623\,
            I => \U712_CHIP_RAM.N_113\
        );

    \I__880\ : CascadeMux
    port map (
            O => \N__5618\,
            I => \N__5614\
        );

    \I__879\ : InMux
    port map (
            O => \N__5617\,
            I => \N__5611\
        );

    \I__878\ : InMux
    port map (
            O => \N__5614\,
            I => \N__5608\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__5611\,
            I => \N__5604\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__5608\,
            I => \N__5601\
        );

    \I__875\ : InMux
    port map (
            O => \N__5607\,
            I => \N__5597\
        );

    \I__874\ : Span4Mux_v
    port map (
            O => \N__5604\,
            I => \N__5592\
        );

    \I__873\ : Span4Mux_v
    port map (
            O => \N__5601\,
            I => \N__5592\
        );

    \I__872\ : InMux
    port map (
            O => \N__5600\,
            I => \N__5589\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__5597\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__870\ : Odrv4
    port map (
            O => \N__5592\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__5589\,
            I => \U712_CHIP_RAM.N_413\
        );

    \I__868\ : IoInMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__866\ : IoSpan4Mux
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__865\ : Sp12to4
    port map (
            O => \N__5573\,
            I => \N__5570\
        );

    \I__864\ : Span12Mux_s7_h
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__863\ : Span12Mux_h
    port map (
            O => \N__5567\,
            I => \N__5563\
        );

    \I__862\ : InMux
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__861\ : Odrv12
    port map (
            O => \N__5563\,
            I => \CLK_EN_c\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__5560\,
            I => \CLK_EN_c\
        );

    \I__859\ : InMux
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__5552\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\
        );

    \I__857\ : CascadeMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__856\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5542\
        );

    \I__855\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__5542\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__853\ : LocalMux
    port map (
            O => \N__5539\,
            I => \U712_CHIP_RAM.N_342\
        );

    \I__852\ : InMux
    port map (
            O => \N__5534\,
            I => \N__5531\
        );

    \I__851\ : LocalMux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__850\ : Odrv4
    port map (
            O => \N__5528\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\
        );

    \I__849\ : InMux
    port map (
            O => \N__5525\,
            I => \N__5521\
        );

    \I__848\ : InMux
    port map (
            O => \N__5524\,
            I => \N__5518\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__5518\,
            I => \N__5512\
        );

    \I__845\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5509\
        );

    \I__844\ : Span4Mux_v
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__843\ : Sp12to4
    port map (
            O => \N__5509\,
            I => \N__5501\
        );

    \I__842\ : Sp12to4
    port map (
            O => \N__5506\,
            I => \N__5501\
        );

    \I__841\ : Span12Mux_h
    port map (
            O => \N__5501\,
            I => \N__5498\
        );

    \I__840\ : Span12Mux_v
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__839\ : Odrv12
    port map (
            O => \N__5495\,
            I => \AWEn_c\
        );

    \I__838\ : IoInMux
    port map (
            O => \N__5492\,
            I => \N__5489\
        );

    \I__837\ : LocalMux
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__836\ : Span4Mux_s3_v
    port map (
            O => \N__5486\,
            I => \N__5483\
        );

    \I__835\ : Span4Mux_v
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__5477\,
            I => \N__5473\
        );

    \I__832\ : InMux
    port map (
            O => \N__5476\,
            I => \N__5470\
        );

    \I__831\ : Odrv4
    port map (
            O => \N__5473\,
            I => \DBDIR_c\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__5470\,
            I => \DBDIR_c\
        );

    \I__829\ : InMux
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__5462\,
            I => \N__5458\
        );

    \I__827\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__826\ : Odrv4
    port map (
            O => \N__5458\,
            I => \DBRn_c_i\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__5455\,
            I => \DBRn_c_i\
        );

    \I__824\ : IoInMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__822\ : Span12Mux_s4_h
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__821\ : Odrv12
    port map (
            O => \N__5441\,
            I => \DBRn_c_i_0\
        );

    \I__820\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5435\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__817\ : Sp12to4
    port map (
            O => \N__5429\,
            I => \N__5426\
        );

    \I__816\ : Odrv12
    port map (
            O => \N__5426\,
            I => \A_c_13\
        );

    \I__815\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__813\ : Span4Mux_v
    port map (
            O => \N__5417\,
            I => \N__5414\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__811\ : Sp12to4
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__810\ : Odrv12
    port map (
            O => \N__5408\,
            I => \A_c_12\
        );

    \I__809\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5402\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__806\ : Span4Mux_v
    port map (
            O => \N__5396\,
            I => \N__5393\
        );

    \I__805\ : Sp12to4
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__804\ : Odrv12
    port map (
            O => \N__5390\,
            I => \A_c_5\
        );

    \I__803\ : InMux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__802\ : LocalMux
    port map (
            O => \N__5384\,
            I => \N__5381\
        );

    \I__801\ : Span4Mux_v
    port map (
            O => \N__5381\,
            I => \N__5378\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__799\ : Sp12to4
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__798\ : Odrv12
    port map (
            O => \N__5372\,
            I => \A_c_15\
        );

    \I__797\ : InMux
    port map (
            O => \N__5369\,
            I => \N__5366\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__5363\,
            I => \N__5360\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__793\ : Sp12to4
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__792\ : Odrv12
    port map (
            O => \N__5354\,
            I => \A_c_8\
        );

    \I__791\ : InMux
    port map (
            O => \N__5351\,
            I => \N__5347\
        );

    \I__790\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__5344\,
            I => \N__5336\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__5341\,
            I => \N__5333\
        );

    \I__786\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5330\
        );

    \I__785\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5327\
        );

    \I__784\ : Odrv4
    port map (
            O => \N__5336\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__783\ : Odrv4
    port map (
            O => \N__5333\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__5330\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__5327\,
            I => \U712_CHIP_RAM.N_261\
        );

    \I__780\ : InMux
    port map (
            O => \N__5318\,
            I => \N__5315\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__5315\,
            I => \N__5312\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__777\ : Sp12to4
    port map (
            O => \N__5309\,
            I => \N__5306\
        );

    \I__776\ : Odrv12
    port map (
            O => \N__5306\,
            I => \A_c_11\
        );

    \I__775\ : InMux
    port map (
            O => \N__5303\,
            I => \N__5300\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5297\
        );

    \I__773\ : Sp12to4
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__772\ : Span12Mux_v
    port map (
            O => \N__5294\,
            I => \N__5291\
        );

    \I__771\ : Span12Mux_h
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__770\ : Odrv12
    port map (
            O => \N__5288\,
            I => \A_c_4\
        );

    \I__769\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5282\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__5282\,
            I => \U712_CHIP_RAM.N_312\
        );

    \I__767\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__5276\,
            I => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0\
        );

    \I__765\ : CascadeMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__764\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__762\ : Span4Mux_h
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__5261\,
            I => \U712_CHIP_RAM.N_314\
        );

    \I__760\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5255\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__5255\,
            I => \N__5251\
        );

    \I__758\ : InMux
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__757\ : Span4Mux_h
    port map (
            O => \N__5251\,
            I => \N__5245\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__5248\,
            I => \U712_CHIP_RAM.N_459\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__5245\,
            I => \U712_CHIP_RAM.N_459\
        );

    \I__754\ : InMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__5237\,
            I => \N__5232\
        );

    \I__752\ : InMux
    port map (
            O => \N__5236\,
            I => \N__5227\
        );

    \I__751\ : InMux
    port map (
            O => \N__5235\,
            I => \N__5227\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__5232\,
            I => \N__5224\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__5227\,
            I => \U712_CHIP_RAM.N_449\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__5224\,
            I => \U712_CHIP_RAM.N_449\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5219\,
            I => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_\
        );

    \I__746\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5211\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__5215\,
            I => \N__5201\
        );

    \I__744\ : InMux
    port map (
            O => \N__5214\,
            I => \N__5197\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__5211\,
            I => \N__5194\
        );

    \I__742\ : InMux
    port map (
            O => \N__5210\,
            I => \N__5189\
        );

    \I__741\ : InMux
    port map (
            O => \N__5209\,
            I => \N__5189\
        );

    \I__740\ : InMux
    port map (
            O => \N__5208\,
            I => \N__5178\
        );

    \I__739\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5178\
        );

    \I__738\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5171\
        );

    \I__737\ : InMux
    port map (
            O => \N__5205\,
            I => \N__5171\
        );

    \I__736\ : InMux
    port map (
            O => \N__5204\,
            I => \N__5171\
        );

    \I__735\ : InMux
    port map (
            O => \N__5201\,
            I => \N__5164\
        );

    \I__734\ : InMux
    port map (
            O => \N__5200\,
            I => \N__5164\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__5197\,
            I => \N__5161\
        );

    \I__732\ : Span4Mux_h
    port map (
            O => \N__5194\,
            I => \N__5156\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__5189\,
            I => \N__5156\
        );

    \I__730\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5153\
        );

    \I__729\ : InMux
    port map (
            O => \N__5187\,
            I => \N__5144\
        );

    \I__728\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5144\
        );

    \I__727\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5144\
        );

    \I__726\ : InMux
    port map (
            O => \N__5184\,
            I => \N__5144\
        );

    \I__725\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5141\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__5178\,
            I => \N__5138\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__5171\,
            I => \N__5135\
        );

    \I__722\ : InMux
    port map (
            O => \N__5170\,
            I => \N__5130\
        );

    \I__721\ : InMux
    port map (
            O => \N__5169\,
            I => \N__5130\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__5164\,
            I => \N__5126\
        );

    \I__719\ : Span4Mux_v
    port map (
            O => \N__5161\,
            I => \N__5121\
        );

    \I__718\ : Span4Mux_v
    port map (
            O => \N__5156\,
            I => \N__5121\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__5153\,
            I => \N__5114\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5114\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5114\
        );

    \I__714\ : Span4Mux_v
    port map (
            O => \N__5138\,
            I => \N__5107\
        );

    \I__713\ : Span4Mux_v
    port map (
            O => \N__5135\,
            I => \N__5107\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__5130\,
            I => \N__5107\
        );

    \I__711\ : InMux
    port map (
            O => \N__5129\,
            I => \N__5104\
        );

    \I__710\ : Span12Mux_v
    port map (
            O => \N__5126\,
            I => \N__5093\
        );

    \I__709\ : Sp12to4
    port map (
            O => \N__5121\,
            I => \N__5093\
        );

    \I__708\ : Span12Mux_v
    port map (
            O => \N__5114\,
            I => \N__5093\
        );

    \I__707\ : Sp12to4
    port map (
            O => \N__5107\,
            I => \N__5093\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__5104\,
            I => \N__5093\
        );

    \I__705\ : Span12Mux_h
    port map (
            O => \N__5093\,
            I => \N__5090\
        );

    \I__704\ : Odrv12
    port map (
            O => \N__5090\,
            I => \RESETn_c\
        );

    \I__703\ : InMux
    port map (
            O => \N__5087\,
            I => \N__5078\
        );

    \I__702\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5078\
        );

    \I__701\ : InMux
    port map (
            O => \N__5085\,
            I => \N__5078\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__5078\,
            I => \N__5074\
        );

    \I__699\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5071\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__5074\,
            I => \U712_CHIP_RAM.N_421\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__5071\,
            I => \U712_CHIP_RAM.N_421\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5066\,
            I => \U712_CYCLE_TERM.N_286_i_0_en_cascade_\
        );

    \I__695\ : IoInMux
    port map (
            O => \N__5063\,
            I => \N__5060\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__693\ : Span12Mux_s1_v
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__692\ : Span12Mux_v
    port map (
            O => \N__5054\,
            I => \N__5050\
        );

    \I__691\ : InMux
    port map (
            O => \N__5053\,
            I => \N__5047\
        );

    \I__690\ : Odrv12
    port map (
            O => \N__5050\,
            I => \RESETn_c_i\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__5047\,
            I => \RESETn_c_i\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5042\,
            I => \N__5038\
        );

    \I__687\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5032\
        );

    \I__686\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5029\
        );

    \I__685\ : InMux
    port map (
            O => \N__5037\,
            I => \N__5022\
        );

    \I__684\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5022\
        );

    \I__683\ : InMux
    port map (
            O => \N__5035\,
            I => \N__5022\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__5032\,
            I => \N__5019\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__5029\,
            I => \N__5016\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__5022\,
            I => \N__5013\
        );

    \I__679\ : Odrv4
    port map (
            O => \N__5019\,
            I => \CPU_TACK\
        );

    \I__678\ : Odrv12
    port map (
            O => \N__5016\,
            I => \CPU_TACK\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__5013\,
            I => \CPU_TACK\
        );

    \I__676\ : CEMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__5003\,
            I => \N__5000\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__5000\,
            I => \U712_CYCLE_TERM.N_286_i_0_en_0\
        );

    \I__673\ : InMux
    port map (
            O => \N__4997\,
            I => \N__4993\
        );

    \I__672\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4989\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__4993\,
            I => \N__4986\
        );

    \I__670\ : InMux
    port map (
            O => \N__4992\,
            I => \N__4983\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__4989\,
            I => \N__4980\
        );

    \I__668\ : Span4Mux_v
    port map (
            O => \N__4986\,
            I => \N__4975\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4975\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__4980\,
            I => \N__4972\
        );

    \I__665\ : Span4Mux_v
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__663\ : Sp12to4
    port map (
            O => \N__4969\,
            I => \N__4963\
        );

    \I__662\ : Sp12to4
    port map (
            O => \N__4966\,
            I => \N__4958\
        );

    \I__661\ : Span12Mux_h
    port map (
            O => \N__4963\,
            I => \N__4958\
        );

    \I__660\ : Odrv12
    port map (
            O => \N__4958\,
            I => \DBRn_c\
        );

    \I__659\ : InMux
    port map (
            O => \N__4955\,
            I => \N__4952\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4952\,
            I => \U712_REG_SM.DBR_SYNCZ0Z_0\
        );

    \I__657\ : InMux
    port map (
            O => \N__4949\,
            I => \N__4946\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4943\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__4943\,
            I => \TACK_EN_i_ess\
        );

    \I__654\ : IoInMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__652\ : IoSpan4Mux
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__651\ : Span4Mux_s3_h
    port map (
            O => \N__4931\,
            I => \N__4928\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__649\ : Span4Mux_h
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__4922\,
            I => \N_977_i\
        );

    \I__647\ : IoInMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__4916\,
            I => \N__4913\
        );

    \I__645\ : Span4Mux_s2_v
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__4910\,
            I => \N__4907\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__4907\,
            I => \N__4904\
        );

    \I__642\ : Odrv4
    port map (
            O => \N__4904\,
            I => \VBENn_c\
        );

    \I__641\ : IoInMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__4898\,
            I => \N__4895\
        );

    \I__639\ : Span4Mux_s2_v
    port map (
            O => \N__4895\,
            I => \N__4892\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__4892\,
            I => \N__4888\
        );

    \I__637\ : InMux
    port map (
            O => \N__4891\,
            I => \N__4885\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__4888\,
            I => \N__4882\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__4885\,
            I => \N__4879\
        );

    \I__634\ : Sp12to4
    port map (
            O => \N__4882\,
            I => \N__4876\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__4879\,
            I => \N__4873\
        );

    \I__632\ : Odrv12
    port map (
            O => \N__4876\,
            I => \CONSTANT_ONE_NET\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__4873\,
            I => \CONSTANT_ONE_NET\
        );

    \I__630\ : InMux
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__628\ : Sp12to4
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__627\ : Span12Mux_v
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__626\ : Span12Mux_h
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__4853\,
            I => \A_c_6\
        );

    \I__624\ : InMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4847\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\
        );

    \I__622\ : InMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__4838\,
            I => \N__4835\
        );

    \I__619\ : Odrv4
    port map (
            O => \N__4835\,
            I => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\
        );

    \I__618\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4828\
        );

    \I__617\ : InMux
    port map (
            O => \N__4831\,
            I => \N__4825\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4828\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4825\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__613\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4814\,
            I => \U712_CYCLE_TERM.TACK_STATE_r_sx_1\
        );

    \I__611\ : InMux
    port map (
            O => \N__4811\,
            I => \N__4806\
        );

    \I__610\ : InMux
    port map (
            O => \N__4810\,
            I => \N__4801\
        );

    \I__609\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4801\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4806\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__4801\,
            I => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\
        );

    \I__606\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4790\
        );

    \I__605\ : InMux
    port map (
            O => \N__4795\,
            I => \N__4790\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4790\,
            I => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4787\,
            I => \U712_CYCLE_TERM.N_286_i_0_0_cascade_\
        );

    \I__602\ : InMux
    port map (
            O => \N__4784\,
            I => \N__4781\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4781\,
            I => \N__4777\
        );

    \I__600\ : InMux
    port map (
            O => \N__4780\,
            I => \N__4773\
        );

    \I__599\ : Span4Mux_v
    port map (
            O => \N__4777\,
            I => \N__4770\
        );

    \I__598\ : InMux
    port map (
            O => \N__4776\,
            I => \N__4767\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__4773\,
            I => \U712_CHIP_RAM.N_416\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__4770\,
            I => \U712_CHIP_RAM.N_416\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__4767\,
            I => \U712_CHIP_RAM.N_416\
        );

    \I__594\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4757\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4757\,
            I => \N__4754\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__4754\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__4751\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_\
        );

    \I__590\ : InMux
    port map (
            O => \N__4748\,
            I => \N__4745\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4745\,
            I => \N__4742\
        );

    \I__588\ : Odrv12
    port map (
            O => \N__4742\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__4739\,
            I => \N__4736\
        );

    \I__586\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4733\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__4733\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0\
        );

    \I__584\ : InMux
    port map (
            O => \N__4730\,
            I => \N__4724\
        );

    \I__583\ : InMux
    port map (
            O => \N__4729\,
            I => \N__4724\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__4724\,
            I => \N__4715\
        );

    \I__581\ : InMux
    port map (
            O => \N__4723\,
            I => \N__4708\
        );

    \I__580\ : InMux
    port map (
            O => \N__4722\,
            I => \N__4708\
        );

    \I__579\ : InMux
    port map (
            O => \N__4721\,
            I => \N__4708\
        );

    \I__578\ : InMux
    port map (
            O => \N__4720\,
            I => \N__4701\
        );

    \I__577\ : InMux
    port map (
            O => \N__4719\,
            I => \N__4701\
        );

    \I__576\ : InMux
    port map (
            O => \N__4718\,
            I => \N__4701\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4715\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4708\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__4701\,
            I => \U712_CHIP_RAM.N_45\
        );

    \I__572\ : CascadeMux
    port map (
            O => \N__4694\,
            I => \U712_CHIP_RAM.N_61_cascade_\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__4691\,
            I => \N__4688\
        );

    \I__570\ : InMux
    port map (
            O => \N__4688\,
            I => \N__4683\
        );

    \I__569\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4680\
        );

    \I__568\ : InMux
    port map (
            O => \N__4686\,
            I => \N__4677\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__4683\,
            I => \N__4674\
        );

    \I__566\ : LocalMux
    port map (
            O => \N__4680\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4677\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__4674\,
            I => \U712_CHIP_RAM.REFRESHZ0\
        );

    \I__563\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__562\ : LocalMux
    port map (
            O => \N__4664\,
            I => \U712_CHIP_RAM.N_263\
        );

    \I__561\ : InMux
    port map (
            O => \N__4661\,
            I => \N__4657\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__4660\,
            I => \N__4653\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4657\,
            I => \N__4650\
        );

    \I__558\ : InMux
    port map (
            O => \N__4656\,
            I => \N__4647\
        );

    \I__557\ : InMux
    port map (
            O => \N__4653\,
            I => \N__4644\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__4650\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4647\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__4644\,
            I => \U712_CHIP_RAM.N_271\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__4637\,
            I => \U712_CHIP_RAM.N_341_cascade_\
        );

    \I__552\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4631\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4631\,
            I => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\
        );

    \I__550\ : InMux
    port map (
            O => \N__4628\,
            I => \N__4625\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__4625\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2\
        );

    \I__548\ : InMux
    port map (
            O => \N__4622\,
            I => \N__4619\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__546\ : Span4Mux_v
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__545\ : Span4Mux_v
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__544\ : Sp12to4
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__543\ : Span12Mux_h
    port map (
            O => \N__4607\,
            I => \N__4604\
        );

    \I__542\ : Odrv12
    port map (
            O => \N__4604\,
            I => \A_c_20\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__4601\,
            I => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\
        );

    \I__540\ : InMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__4595\,
            I => \U712_CHIP_RAM.N_362\
        );

    \I__538\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4588\
        );

    \I__537\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4585\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__4588\,
            I => \U712_CHIP_RAM.N_470\
        );

    \I__535\ : LocalMux
    port map (
            O => \N__4585\,
            I => \U712_CHIP_RAM.N_470\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__4580\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_\
        );

    \I__533\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__4574\,
            I => \U712_CHIP_RAM.N_344\
        );

    \I__531\ : InMux
    port map (
            O => \N__4571\,
            I => \N__4568\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4568\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__4565\,
            I => \U712_CHIP_RAM.N_344_cascade_\
        );

    \I__528\ : CascadeMux
    port map (
            O => \N__4562\,
            I => \N__4558\
        );

    \I__527\ : InMux
    port map (
            O => \N__4561\,
            I => \N__4554\
        );

    \I__526\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4551\
        );

    \I__525\ : InMux
    port map (
            O => \N__4557\,
            I => \N__4548\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__4554\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4551\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__522\ : LocalMux
    port map (
            O => \N__4548\,
            I => \U712_CHIP_RAM.N_267\
        );

    \I__521\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4538\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__4535\,
            I => \U712_CHIP_RAM.N_333\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__4532\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_\
        );

    \I__517\ : InMux
    port map (
            O => \N__4529\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\
        );

    \I__516\ : InMux
    port map (
            O => \N__4526\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\
        );

    \I__515\ : InMux
    port map (
            O => \N__4523\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\
        );

    \I__514\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4516\
        );

    \I__513\ : InMux
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__4516\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__4513\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\
        );

    \I__510\ : InMux
    port map (
            O => \N__4508\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\
        );

    \I__509\ : InMux
    port map (
            O => \N__4505\,
            I => \N__4501\
        );

    \I__508\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4498\
        );

    \I__507\ : LocalMux
    port map (
            O => \N__4501\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__4498\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\
        );

    \I__505\ : InMux
    port map (
            O => \N__4493\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\
        );

    \I__504\ : InMux
    port map (
            O => \N__4490\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\
        );

    \I__503\ : InMux
    port map (
            O => \N__4487\,
            I => \N__4483\
        );

    \I__502\ : InMux
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__501\ : LocalMux
    port map (
            O => \N__4483\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__4480\,
            I => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\
        );

    \I__499\ : IoInMux
    port map (
            O => \N__4475\,
            I => \N__4472\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__497\ : Span4Mux_s2_v
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__496\ : Sp12to4
    port map (
            O => \N__4466\,
            I => \N__4463\
        );

    \I__495\ : Span12Mux_h
    port map (
            O => \N__4463\,
            I => \N__4460\
        );

    \I__494\ : Odrv12
    port map (
            O => \N__4460\,
            I => \BANK0_c\
        );

    \I__493\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4453\
        );

    \I__492\ : InMux
    port map (
            O => \N__4456\,
            I => \N__4450\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__4453\,
            I => \U712_CHIP_RAM.N_404\
        );

    \I__490\ : LocalMux
    port map (
            O => \N__4450\,
            I => \U712_CHIP_RAM.N_404\
        );

    \I__489\ : CascadeMux
    port map (
            O => \N__4445\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\
        );

    \I__488\ : InMux
    port map (
            O => \N__4442\,
            I => \N__4438\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__4441\,
            I => \N__4435\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__4438\,
            I => \N__4432\
        );

    \I__485\ : InMux
    port map (
            O => \N__4435\,
            I => \N__4429\
        );

    \I__484\ : Odrv12
    port map (
            O => \N__4432\,
            I => \LATCH_RAM\
        );

    \I__483\ : LocalMux
    port map (
            O => \N__4429\,
            I => \LATCH_RAM\
        );

    \I__482\ : IoInMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__480\ : Span12Mux_s11_v
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__479\ : Odrv12
    port map (
            O => \N__4415\,
            I => \LATCH_CLK_0_i\
        );

    \I__478\ : CascadeMux
    port map (
            O => \N__4412\,
            I => \U712_CHIP_RAM.N_296_cascade_\
        );

    \I__477\ : InMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__4406\,
            I => \U712_CHIP_RAM.N_296\
        );

    \I__475\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__474\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__473\ : Span4Mux_v
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__472\ : Odrv4
    port map (
            O => \N__4394\,
            I => \U712_CHIP_RAM.N_63\
        );

    \I__471\ : InMux
    port map (
            O => \N__4391\,
            I => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\
        );

    \I__470\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4383\
        );

    \I__469\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4378\
        );

    \I__468\ : InMux
    port map (
            O => \N__4386\,
            I => \N__4378\
        );

    \I__467\ : LocalMux
    port map (
            O => \N__4383\,
            I => \N__4375\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__4378\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__465\ : Odrv4
    port map (
            O => \N__4375\,
            I => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\
        );

    \I__464\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__4367\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\
        );

    \I__462\ : IoInMux
    port map (
            O => \N__4364\,
            I => \N__4361\
        );

    \I__461\ : LocalMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__460\ : IoSpan4Mux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__458\ : Span12Mux_s6_h
    port map (
            O => \N__4352\,
            I => \N__4349\
        );

    \I__457\ : Span12Mux_v
    port map (
            O => \N__4349\,
            I => \N__4345\
        );

    \I__456\ : InMux
    port map (
            O => \N__4348\,
            I => \N__4342\
        );

    \I__455\ : Odrv12
    port map (
            O => \N__4345\,
            I => \TACK_OUTn\
        );

    \I__454\ : LocalMux
    port map (
            O => \N__4342\,
            I => \TACK_OUTn\
        );

    \I__453\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__4334\,
            I => \DBR_SYNCZ0Z_0\
        );

    \I__451\ : InMux
    port map (
            O => \N__4331\,
            I => \N__4327\
        );

    \I__450\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4324\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__4327\,
            I => \N__4321\
        );

    \I__448\ : LocalMux
    port map (
            O => \N__4324\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__447\ : Odrv12
    port map (
            O => \N__4321\,
            I => \DBR_SYNCZ0Z_1\
        );

    \I__446\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4311\
        );

    \I__445\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4308\
        );

    \I__444\ : IoInMux
    port map (
            O => \N__4314\,
            I => \N__4305\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__4311\,
            I => \N__4300\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__4308\,
            I => \N__4300\
        );

    \I__441\ : LocalMux
    port map (
            O => \N__4305\,
            I => \N__4297\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__4300\,
            I => \N__4294\
        );

    \I__439\ : Span12Mux_s3_h
    port map (
            O => \N__4297\,
            I => \N__4291\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__4294\,
            I => \N__4288\
        );

    \I__437\ : Span12Mux_v
    port map (
            O => \N__4291\,
            I => \N__4285\
        );

    \I__436\ : Span12Mux_h
    port map (
            O => \N__4288\,
            I => \N__4282\
        );

    \I__435\ : Span12Mux_h
    port map (
            O => \N__4285\,
            I => \N__4279\
        );

    \I__434\ : Span12Mux_v
    port map (
            O => \N__4282\,
            I => \N__4276\
        );

    \I__433\ : Odrv12
    port map (
            O => \N__4279\,
            I => \CLK40_PLL\
        );

    \I__432\ : Odrv12
    port map (
            O => \N__4276\,
            I => \CLK40_PLL\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__430\ : InMux
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__4265\,
            I => \N__4262\
        );

    \I__428\ : Odrv12
    port map (
            O => \N__4262\,
            I => \U712_BYTE_ENABLE.N_90\
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__4259\,
            I => \N__4255\
        );

    \I__426\ : InMux
    port map (
            O => \N__4258\,
            I => \N__4250\
        );

    \I__425\ : InMux
    port map (
            O => \N__4255\,
            I => \N__4250\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__4250\,
            I => \N__4240\
        );

    \I__423\ : ClkMux
    port map (
            O => \N__4249\,
            I => \N__4223\
        );

    \I__422\ : ClkMux
    port map (
            O => \N__4248\,
            I => \N__4223\
        );

    \I__421\ : ClkMux
    port map (
            O => \N__4247\,
            I => \N__4223\
        );

    \I__420\ : ClkMux
    port map (
            O => \N__4246\,
            I => \N__4223\
        );

    \I__419\ : ClkMux
    port map (
            O => \N__4245\,
            I => \N__4223\
        );

    \I__418\ : ClkMux
    port map (
            O => \N__4244\,
            I => \N__4223\
        );

    \I__417\ : ClkMux
    port map (
            O => \N__4243\,
            I => \N__4223\
        );

    \I__416\ : Glb2LocalMux
    port map (
            O => \N__4240\,
            I => \N__4223\
        );

    \I__415\ : GlobalMux
    port map (
            O => \N__4223\,
            I => \N__4220\
        );

    \I__414\ : gio2CtrlBuf
    port map (
            O => \N__4220\,
            I => \CLK40_PLL_g\
        );

    \I__413\ : IoInMux
    port map (
            O => \N__4217\,
            I => \N__4213\
        );

    \I__412\ : IoInMux
    port map (
            O => \N__4216\,
            I => \N__4210\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4205\
        );

    \I__410\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4205\
        );

    \I__409\ : IoSpan4Mux
    port map (
            O => \N__4205\,
            I => \N__4201\
        );

    \I__408\ : IoInMux
    port map (
            O => \N__4204\,
            I => \N__4198\
        );

    \I__407\ : Span4Mux_s2_v
    port map (
            O => \N__4201\,
            I => \N__4195\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__4198\,
            I => \N__4192\
        );

    \I__405\ : Sp12to4
    port map (
            O => \N__4195\,
            I => \N__4189\
        );

    \I__404\ : IoSpan4Mux
    port map (
            O => \N__4192\,
            I => \N__4186\
        );

    \I__403\ : Span12Mux_v
    port map (
            O => \N__4189\,
            I => \N__4183\
        );

    \I__402\ : Span4Mux_s3_h
    port map (
            O => \N__4186\,
            I => \N__4180\
        );

    \I__401\ : Span12Mux_h
    port map (
            O => \N__4183\,
            I => \N__4177\
        );

    \I__400\ : Span4Mux_h
    port map (
            O => \N__4180\,
            I => \N__4174\
        );

    \I__399\ : Odrv12
    port map (
            O => \N__4177\,
            I => \CLK40_PLL_iso_i\
        );

    \I__398\ : Odrv4
    port map (
            O => \N__4174\,
            I => \CLK40_PLL_iso_i\
        );

    \I__397\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__4166\,
            I => \U712_CHIP_RAM.N_414\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__4163\,
            I => \U712_CHIP_RAM.N_415_cascade_\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__4160\,
            I => \U712_CHIP_RAM.N_373_cascade_\
        );

    \I__393\ : CascadeMux
    port map (
            O => \N__4157\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\
        );

    \I__392\ : CEMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__4151\,
            I => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\
        );

    \I__390\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__389\ : LocalMux
    port map (
            O => \N__4145\,
            I => \U712_CHIP_RAM.N_373\
        );

    \I__388\ : IoInMux
    port map (
            O => \N__4142\,
            I => \N__4139\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__386\ : IoSpan4Mux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__385\ : Span4Mux_s2_v
    port map (
            O => \N__4133\,
            I => \N__4130\
        );

    \I__384\ : Sp12to4
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__383\ : Odrv12
    port map (
            O => \N__4127\,
            I => \N_48_i\
        );

    \I__382\ : InMux
    port map (
            O => \N__4124\,
            I => \N__4121\
        );

    \I__381\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4118\
        );

    \I__380\ : Span12Mux_v
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__379\ : Odrv12
    port map (
            O => \N__4115\,
            I => \RAMSPACEn_c\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__4112\,
            I => \U712_CHIP_RAM.N_355_cascade_\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__4109\,
            I => \U712_CHIP_RAM.N_416_cascade_\
        );

    \I__376\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__4103\,
            I => \U712_CHIP_RAM.N_448\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__4100\,
            I => \U712_CHIP_RAM.N_261_cascade_\
        );

    \I__373\ : CascadeMux
    port map (
            O => \N__4097\,
            I => \U712_CHIP_RAM.N_404_cascade_\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__4094\,
            I => \U712_CHIP_RAM.N_413_cascade_\
        );

    \I__371\ : IoInMux
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__369\ : Span4Mux_s2_v
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__368\ : Span4Mux_v
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__4079\,
            I => \CLK80_PLL_i_i\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__4076\,
            I => \U712_CHIP_RAM.N_448_cascade_\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__4073\,
            I => \U712_CHIP_RAM.N_459_cascade_\
        );

    \I__364\ : CascadeMux
    port map (
            O => \N__4070\,
            I => \U712_CHIP_RAM.N_308_cascade_\
        );

    \I__363\ : InMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__4064\,
            I => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\
        );

    \I__361\ : IoInMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__359\ : Span4Mux_s0_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__358\ : Span4Mux_v
    port map (
            O => \N__4052\,
            I => \N__4049\
        );

    \I__357\ : Sp12to4
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__356\ : Span12Mux_h
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__355\ : Span12Mux_v
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__354\ : Odrv12
    port map (
            O => \N__4040\,
            I => \CLK40_IN_c\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            I => \N__7673\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            I => \N__7675\
        );

    \INVU712_REG_SM.REG_CYCLE_STARTC\ : INV
    port map (
            O => \INVU712_REG_SM.REG_CYCLE_STARTC_net\,
            I => \N__4244\
        );

    \INVU712_REG_SM.UDSnC\ : INV
    port map (
            O => \INVU712_REG_SM.UDSnC_net\,
            I => \N__4243\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            I => \N__7676\
        );

    \INVU712_REG_SM.C3_SYNC_0C\ : INV
    port map (
            O => \INVU712_REG_SM.C3_SYNC_0C_net\,
            I => \N__4245\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            I => \N__7677\
        );

    \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            I => \N__7679\
        );

    \INVU712_REG_SM.STATE_COUNTER_2C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            I => \N__4248\
        );

    \INVU712_REG_SM.REG_CYCLEC\ : INV
    port map (
            O => \INVU712_REG_SM.REG_CYCLEC_net\,
            I => \N__4247\
        );

    \INVU712_REG_SM.STATE_COUNTER_5C\ : INV
    port map (
            O => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            I => \N__4246\
        );

    \INVU712_CHIP_RAM.DMA_A20C\ : INV
    port map (
            O => \INVU712_CHIP_RAM.DMA_A20C_net\,
            I => \N__7678\
        );

    \INVU712_REG_SM.DBR_SYNC_1C\ : INV
    port map (
            O => \INVU712_REG_SM.DBR_SYNC_1C_net\,
            I => \N__4249\
        );

    \IN_MUX_bfv_12_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_10_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_8_0_\
        );

    \C1_ibuf_RNIPA2A\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7516\,
            GLOBALBUFFEROUTPUT => \C1_c_g\
        );

    \CLK40_PLL_derived_clock_RNIIOT\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__4314\,
            GLOBALBUFFEROUTPUT => \CLK40_PLL_g\
        );

    \RESETn_ibuf_RNIM9SF_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5063\,
            GLOBALBUFFEROUTPUT => \RESETn_c_i_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \DBRn_c_i_0_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__5450\,
            GLOBALBUFFEROUTPUT => \DBRn_c_i_0_g\
        );

    \C3_ibuf_RNIRKME\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__7151\,
            GLOBALBUFFEROUTPUT => \C3_c_g\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \CLKRAM_obuf_RNO_LC_3_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__9743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK80_PLL_i_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBR_SYNC_0_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4996\,
            lcout => \DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9737\,
            ce => 'H',
            sr => \N__10992\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_1_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101010110101"
        )
    port map (
            in0 => \N__6473\,
            in1 => \N__6626\,
            in2 => \N__6406\,
            in3 => \N__6192\,
            lcout => \U712_CHIP_RAM.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__6193\,
            in1 => \N__4780\,
            in2 => \N__6293\,
            in3 => \N__6096\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI8UIP2_4_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__6471\,
            in1 => \N__6687\,
            in2 => \N__5907\,
            in3 => \N__5339\,
            lcout => \U712_CHIP_RAM.N_448\,
            ltout => \U712_CHIP_RAM.N_448_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI4CEN3_0_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6617\,
            in2 => \N__4076\,
            in3 => \N__6388\,
            lcout => \U712_CHIP_RAM.N_459\,
            ltout => \U712_CHIP_RAM.N_459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010100000"
        )
    port map (
            in0 => \N__5207\,
            in1 => \_gnd_net_\,
            in2 => \N__4073\,
            in3 => \N__6200\,
            lcout => \U712_CHIP_RAM.SDRAM_CONFIGUREDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNO_0_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__6267\,
            in1 => \N__5525\,
            in2 => \_gnd_net_\,
            in3 => \N__7934\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_308_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_LC_7_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__5208\,
            in1 => \N__7410\,
            in2 => \N__4070\,
            in3 => \N__4067\,
            lcout => \WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9726\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNIEH9V_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__4331\,
            in1 => \N__4686\,
            in2 => \_gnd_net_\,
            in3 => \N__4388\,
            lcout => \U712_CHIP_RAM.N_416\,
            ltout => \U712_CHIP_RAM.N_416_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6266\,
            in2 => \N__4109\,
            in3 => \N__4656\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_8_i_i_a3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNISAAQ_4_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5891\,
            in2 => \_gnd_net_\,
            in3 => \N__6160\,
            lcout => \U712_CHIP_RAM.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIJIDU3_0_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6360\,
            in1 => \N__4106\,
            in2 => \N__4562\,
            in3 => \N__10635\,
            lcout => \U712_CHIP_RAM.N_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI94JE1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7000\,
            in1 => \N__6571\,
            in2 => \N__6719\,
            in3 => \N__5893\,
            lcout => \U712_CHIP_RAM.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI9KPC1_7_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4486\,
            in1 => \N__4504\,
            in2 => \_gnd_net_\,
            in3 => \N__4519\,
            lcout => \U712_CHIP_RAM.N_261\,
            ltout => \U712_CHIP_RAM.N_261_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI41LA2_1_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6445\,
            in2 => \N__4100\,
            in3 => \N__6358\,
            lcout => \U712_CHIP_RAM.N_404\,
            ltout => \U712_CHIP_RAM.N_404_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI0CV43_4_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__5892\,
            in1 => \_gnd_net_\,
            in2 => \N__4097\,
            in3 => \N__6161\,
            lcout => \U712_CHIP_RAM.N_449\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3FV43_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__6688\,
            in1 => \N__5340\,
            in2 => \N__4660\,
            in3 => \N__6446\,
            lcout => \U712_CHIP_RAM.N_413\,
            ltout => \U712_CHIP_RAM.N_413_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIPJCN3_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__6359\,
            in1 => \_gnd_net_\,
            in2 => \N__4094\,
            in3 => \N__7406\,
            lcout => \U712_CHIP_RAM.N_470\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIC9HD1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__6720\,
            in1 => \N__6294\,
            in2 => \_gnd_net_\,
            in3 => \N__6581\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CONFIGURED_RNIKV5I5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__6202\,
            in1 => \N__4169\,
            in2 => \N__4163\,
            in3 => \N__4457\,
            lcout => \U712_CHIP_RAM.N_373\,
            ltout => \U712_CHIP_RAM.N_373_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNICBGO9_2_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6582\,
            in2 => \N__4160\,
            in3 => \N__4591\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0\,
            ltout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNO_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4157\,
            in3 => \N__11029\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_10_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6093\,
            in1 => \N__6203\,
            in2 => \_gnd_net_\,
            in3 => \N__6295\,
            lcout => \DMA_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9730\,
            ce => \N__4154\,
            sr => \N__11000\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_1_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101010101010"
        )
    port map (
            in0 => \N__4148\,
            in1 => \N__4561\,
            in2 => \N__6404\,
            in3 => \N__5607\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_48_i_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100110001011111"
        )
    port map (
            in0 => \N__10646\,
            in1 => \N__10784\,
            in2 => \N__4271\,
            in3 => \N__6943\,
            lcout => \N_48_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNO_0_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__4387\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10645\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_355_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__4124\,
            in1 => \N__5169\,
            in2 => \N__4112\,
            in3 => \N__8011\,
            lcout => \U712_CHIP_RAM.CPU_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_CYCLE_START_RNI0N9G_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4330\,
            in2 => \_gnd_net_\,
            in3 => \N__4386\,
            lcout => \U712_CHIP_RAM.N_263\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_RAM_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010100000"
        )
    port map (
            in0 => \N__5170\,
            in1 => \N__4403\,
            in2 => \N__4441\,
            in3 => \N__4370\,
            lcout => \LATCH_RAM\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9732\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_OUTn_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111110001010"
        )
    port map (
            in0 => \N__4348\,
            in1 => \N__4315\,
            in2 => \N__5840\,
            in3 => \N__4811\,
            lcout => \TACK_OUTn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9735\,
            ce => 'H',
            sr => \N__10987\
        );

    \DBR_SYNC_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4337\,
            lcout => \DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9735\,
            ce => 'H',
            sr => \N__10987\
        );

    \U712_CYCLE_TERM.TACK_STATE_3_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5205\,
            in2 => \_gnd_net_\,
            in3 => \N__4832\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101110111"
        )
    port map (
            in0 => \N__5206\,
            in1 => \N__5789\,
            in2 => \N__4259\,
            in3 => \N__5833\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_r_sx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_2_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5204\,
            in1 => \N__4316\,
            in2 => \_gnd_net_\,
            in3 => \N__5834\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9738\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LLBE_i_o4_0_o3_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110111100101"
        )
    port map (
            in0 => \N__10244\,
            in1 => \N__10319\,
            in2 => \N__10424\,
            in3 => \N__10141\,
            lcout => \U712_BYTE_ENABLE.N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK40_PLL_derived_clock_RNIIOT_0_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__4258\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CLK40_PLL_iso_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.LATCH_CLK_0_i_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5762\,
            in2 => \_gnd_net_\,
            in3 => \N__4442\,
            lcout => \LATCH_CLK_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__7697\,
            in1 => \N__7547\,
            in2 => \N__5215\,
            in3 => \N__6956\,
            lcout => \U712_CHIP_RAM.REFRESHZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111010101010"
        )
    port map (
            in0 => \N__6269\,
            in1 => \N__4844\,
            in2 => \N__7013\,
            in3 => \N__5200\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9723\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_1_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101100000"
        )
    port map (
            in0 => \N__6195\,
            in1 => \N__6475\,
            in2 => \N__6629\,
            in3 => \N__6739\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_1_63_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIRILU_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4687\,
            in2 => \_gnd_net_\,
            in3 => \N__6268\,
            lcout => \U712_CHIP_RAM.N_296\,
            ltout => \U712_CHIP_RAM.N_296_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_1_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011001100"
        )
    port map (
            in0 => \N__6474\,
            in1 => \N__5904\,
            in2 => \N__4412\,
            in3 => \N__6196\,
            lcout => \U712_CHIP_RAM.N_312\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_0_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__4409\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6194\,
            lcout => \U712_CHIP_RAM.N_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.LATCH_RAM_RNO_0_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6389\,
            in2 => \_gnd_net_\,
            in3 => \N__7001\,
            lcout => \U712_CHIP_RAM.N_63\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_1_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6472\,
            in2 => \_gnd_net_\,
            in3 => \N__4391\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_0_2_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6613\,
            in2 => \_gnd_net_\,
            in3 => \N__4529\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER_s_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_3_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4718\,
            in1 => \N__6736\,
            in2 => \_gnd_net_\,
            in3 => \N__4526\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            clk => \N__9725\,
            ce => \N__5680\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_4_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4729\,
            in1 => \N__5906\,
            in2 => \_gnd_net_\,
            in3 => \N__4523\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            clk => \N__9725\,
            ce => \N__5680\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_5_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4719\,
            in1 => \N__4520\,
            in2 => \_gnd_net_\,
            in3 => \N__4508\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            clk => \N__9725\,
            ce => \N__5680\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_6_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4730\,
            in1 => \N__4505\,
            in2 => \_gnd_net_\,
            in3 => \N__4493\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.SDRAM_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.SDRAM_COUNTER_cry_6\,
            clk => \N__9725\,
            ce => \N__5680\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_7_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__4720\,
            in1 => \N__4487\,
            in2 => \_gnd_net_\,
            in3 => \N__4490\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9725\,
            ce => \N__5680\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__4598\,
            in1 => \N__6297\,
            in2 => \N__6095\,
            in3 => \N__5662\,
            lcout => \BANK0_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9727\,
            ce => \N__5645\,
            sr => \N__11001\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI3IG83_3_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__6692\,
            in1 => \_gnd_net_\,
            in2 => \N__6606\,
            in3 => \N__4456\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTER15\,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIURFN4_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4776\,
            in2 => \N__4445\,
            in3 => \N__6296\,
            lcout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa\,
            ltout => \U712_CHIP_RAM.WRITE_CYCLE_2_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__4622\,
            in1 => \_gnd_net_\,
            in2 => \N__4601\,
            in3 => \N__9971\,
            lcout => \U712_CHIP_RAM.N_362\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0AC7_3_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000010"
        )
    port map (
            in0 => \N__5214\,
            in1 => \N__5236\,
            in2 => \N__6094\,
            in3 => \N__6694\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_1_sqmuxa_1_i_0_i_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIUMPVI_3_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__5254\,
            in1 => \N__4592\,
            in2 => \N__4580\,
            in3 => \N__4577\,
            lcout => \U712_CHIP_RAM.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_esr_RNI8MK44_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6987\,
            in1 => \N__6693\,
            in2 => \N__6627\,
            in3 => \N__5235\,
            lcout => \U712_CHIP_RAM.N_344\,
            ltout => \U712_CHIP_RAM.N_344_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__4571\,
            in1 => \N__5545\,
            in2 => \N__4565\,
            in3 => \N__6077\,
            lcout => \U712_CHIP_RAM.N_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIOBA64_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4557\,
            in1 => \N__6370\,
            in2 => \_gnd_net_\,
            in3 => \N__5600\,
            lcout => \U712_CHIP_RAM.N_342\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.WRITE_CYCLE_RNIO6DI_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7416\,
            in2 => \_gnd_net_\,
            in3 => \N__6567\,
            lcout => \U712_CHIP_RAM.N_267\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNO_1_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4891\,
            in2 => \_gnd_net_\,
            in3 => \N__6371\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_COUNTER_s_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__5087\,
            in1 => \N__4541\,
            in2 => \N__4532\,
            in3 => \N__4721\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9729\,
            ce => \N__5684\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIMQBQ1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__4784\,
            in1 => \N__6298\,
            in2 => \_gnd_net_\,
            in3 => \N__6207\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_0_sqmuxa_1_0_a2_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_1_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5085\,
            in1 => \N__4760\,
            in2 => \N__4751\,
            in3 => \N__4722\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9729\,
            ce => \N__5684\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_2_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__5086\,
            in1 => \N__4748\,
            in2 => \N__4739\,
            in3 => \N__4723\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9729\,
            ce => \N__5684\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_1_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__7418\,
            in1 => \N__10573\,
            in2 => \N__6740\,
            in3 => \N__5638\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_61_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011000000"
        )
    port map (
            in0 => \N__5041\,
            in1 => \N__5129\,
            in2 => \N__4694\,
            in3 => \N__4634\,
            lcout => \CPU_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9731\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNIMQBQ1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__6276\,
            in1 => \N__6201\,
            in2 => \N__4691\,
            in3 => \N__4667\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_0_a3_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_2_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6730\,
            in1 => \N__7417\,
            in2 => \_gnd_net_\,
            in3 => \N__6373\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4628\,
            in1 => \N__4661\,
            in2 => \N__4637\,
            in3 => \N__5350\,
            lcout => \U712_CHIP_RAM.CPU_TACK_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CPU_TACK_RNO_3_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111001111111"
        )
    port map (
            in0 => \N__6372\,
            in1 => \N__6599\,
            in2 => \N__6489\,
            in3 => \N__6729\,
            lcout => \U712_CHIP_RAM.un1_SDRAM_COUNTER48_2_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DBRn_ibuf_RNIBAB_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4997\,
            lcout => \DBRn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_1_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4796\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5183\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9733\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNO_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4850\,
            in2 => \_gnd_net_\,
            in3 => \N__4795\,
            lcout => \U712_CHIP_RAM.DMA_CYCLE_START_RNOZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_RNO_0_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4831\,
            in1 => \N__5036\,
            in2 => \N__5839\,
            in3 => \N__4809\,
            lcout => \U712_CYCLE_TERM.TACK_STATE_srsts_0_i_a3_0_1_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001110"
        )
    port map (
            in0 => \N__5037\,
            in1 => \N__6879\,
            in2 => \N__4820\,
            in3 => \N__5832\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_4_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5187\,
            in2 => \_gnd_net_\,
            in3 => \N__4810\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CAS_SYNC_0_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__5185\,
            in1 => \N__10783\,
            in2 => \_gnd_net_\,
            in3 => \N__10868\,
            lcout => \U712_CHIP_RAM.CAS_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9736\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RESETn_ibuf_RNIM9SF_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5184\,
            lcout => \RESETn_c_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_2_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5784\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_286_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_1_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__5800\,
            in1 => \N__5035\,
            in2 => \N__4787\,
            in3 => \N__6878\,
            lcout => OPEN,
            ltout => \U712_CYCLE_TERM.N_286_i_0_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_RNO_0_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5066\,
            in3 => \N__5053\,
            lcout => \U712_CYCLE_TERM.N_286_i_0_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_EN_i_ess_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0111011101111111"
        )
    port map (
            in0 => \N__5188\,
            in1 => \N__5788\,
            in2 => \N__5042\,
            in3 => \N__6881\,
            lcout => \TACK_EN_i_ess\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9739\,
            ce => \N__5006\,
            sr => \N__10979\
        );

    \U712_REG_SM.DBR_SYNC_1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4955\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.DBR_SYNC_1C_net\,
            ce => 'H',
            sr => \N__10977\
        );

    \U712_REG_SM.DBR_SYNC_0_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__4992\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.DBR_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.DBR_SYNC_1C_net\,
            ce => 'H',
            sr => \N__10977\
        );

    \TACKn_obuft_RNO_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4949\,
            lcout => \N_977_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.un1_VBENn_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__10690\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5744\,
            lcout => \VBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIRUMR1_4_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__6622\,
            in1 => \N__6403\,
            in2 => \N__6497\,
            in3 => \N__5905\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_o3_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_4_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4868\,
            in1 => \N__5438\,
            in2 => \_gnd_net_\,
            in3 => \N__9040\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_3_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9037\,
            in1 => \N__5423\,
            in2 => \_gnd_net_\,
            in3 => \N__5405\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_6_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5387\,
            in1 => \N__5369\,
            in2 => \_gnd_net_\,
            in3 => \N__9039\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIVTLS1_7_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5216\,
            in2 => \_gnd_net_\,
            in3 => \N__5351\,
            lcout => \U712_CHIP_RAM.N_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_2_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5318\,
            in1 => \N__5303\,
            in2 => \_gnd_net_\,
            in3 => \N__9038\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_1_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5285\,
            in1 => \N__5279\,
            in2 => \N__5273\,
            in3 => \N__5954\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9724\,
            ce => \N__5935\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNI6VAGA_2_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__5258\,
            in1 => \N__6618\,
            in2 => \N__5618\,
            in3 => \N__5240\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIBVVIG_2_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__5699\,
            in1 => \N__5209\,
            in2 => \N__5219\,
            in3 => \N__5077\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_3_sqmuxa_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPRCO3_3_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5210\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6076\,
            lcout => \U712_CHIP_RAM.N_421\,
            ltout => \U712_CHIP_RAM.N_421_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIB13D6_4_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100011111"
        )
    port map (
            in0 => \N__5698\,
            in1 => \N__5900\,
            in2 => \N__5687\,
            in3 => \N__6212\,
            lcout => \U712_CHIP_RAM.SDRAM_COUNTERe_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_A20_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__9970\,
            in1 => \N__5465\,
            in2 => \N__9413\,
            in3 => \N__5663\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_A20C_net\,
            ce => 'H',
            sr => \N__10993\
        );

    \U712_CHIP_RAM.BANK0_esr_RNO_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11028\,
            in2 => \_gnd_net_\,
            in3 => \N__5651\,
            lcout => \U712_CHIP_RAM.N_18_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CLK_EN_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100010111001100"
        )
    port map (
            in0 => \N__5639\,
            in1 => \N__5566\,
            in2 => \N__6405\,
            in3 => \N__5617\,
            lcout => \CLK_EN_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9728\,
            ce => 'H',
            sr => \N__10988\
        );

    \U712_CHIP_RAM.CPU_CYCLE_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010101100"
        )
    port map (
            in0 => \N__5555\,
            in1 => \N__10574\,
            in2 => \N__5549\,
            in3 => \N__6224\,
            lcout => \CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9728\,
            ce => 'H',
            sr => \N__10988\
        );

    \U712_CHIP_RAM.DBENn_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0100111011101110"
        )
    port map (
            in0 => \N__5534\,
            in1 => \N__7031\,
            in2 => \N__6101\,
            in3 => \N__8501\,
            lcout => \DBENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9728\,
            ce => 'H',
            sr => \N__10988\
        );

    \U712_CHIP_RAM.DBDIR_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__5524\,
            in1 => \N__5476\,
            in2 => \_gnd_net_\,
            in3 => \N__6041\,
            lcout => \DBDIR_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9728\,
            ce => 'H',
            sr => \N__10988\
        );

    \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__7032\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7012\,
            lcout => \U712_BYTE_ENABLE.un1_CLLBEn_i_0_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_ctle_9_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5461\,
            lcout => \DBRn_c_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CYCLE_TERM.TACK_STATE_0_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "0011000010111010"
        )
    port map (
            in0 => \N__5846\,
            in1 => \N__5835\,
            in2 => \N__5804\,
            in3 => \N__6880\,
            lcout => \U712_CYCLE_TERM.TACK_STATEZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9734\,
            ce => 'H',
            sr => \N__10980\
        );

    \U712_REG_SM.STATE_COUNTER_5_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__6800\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10978\
        );

    \U712_REG_SM.STATE_COUNTER_6_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5768\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10978\
        );

    \U712_REG_SM.LATCH_REG_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__5755\,
            in1 => \N__7880\,
            in2 => \N__6785\,
            in3 => \N__8087\,
            lcout => \LATCH_REG\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10978\
        );

    \U712_REG_SM.REG_CPU_CYCLE_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111000000101"
        )
    port map (
            in0 => \N__6799\,
            in1 => \N__5737\,
            in2 => \N__7214\,
            in3 => \N__5723\,
            lcout => \REG_CPU_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_5C_net\,
            ce => 'H',
            sr => \N__10978\
        );

    \U712_REG_SM.DBR_SYNC_RNIVIGC1_1_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__8376\,
            in1 => \N__6753\,
            in2 => \N__8332\,
            in3 => \N__8255\,
            lcout => \U712_REG_SM.STATE_COUNTERc_0\,
            ltout => \U712_REG_SM.STATE_COUNTERc_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CPU_CYCLE_RNO_0_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000111"
        )
    port map (
            in0 => \N__7875\,
            in1 => \N__6798\,
            in2 => \N__5726\,
            in3 => \N__8076\,
            lcout => \U712_REG_SM.REG_CPU_CYCLE_e_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_0_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8377\,
            in1 => \N__6834\,
            in2 => \_gnd_net_\,
            in3 => \N__7874\,
            lcout => \U712_REG_SM.N_297\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_1_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5717\,
            in1 => \N__6035\,
            in2 => \_gnd_net_\,
            in3 => \N__9075\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIMUKI_0_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__9171\,
            in1 => \N__8914\,
            in2 => \_gnd_net_\,
            in3 => \N__9067\,
            lcout => \U712_CHIP_RAM.CMA_5_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_7_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__6020\,
            in1 => \N__6005\,
            in2 => \_gnd_net_\,
            in3 => \N__9066\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_3_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__9068\,
            in1 => \N__5990\,
            in2 => \N__10674\,
            in3 => \N__7067\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_0_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6305\,
            in1 => \N__6641\,
            in2 => \N__5974\,
            in3 => \N__5951\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9719\,
            ce => \N__5936\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_3_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6503\,
            in1 => \N__5981\,
            in2 => \N__5975\,
            in3 => \N__5953\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9719\,
            ce => \N__5936\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIP0891_1_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__6737\,
            in1 => \N__6490\,
            in2 => \_gnd_net_\,
            in3 => \N__6221\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_411_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_COUNTER_RNIPB1M2_4_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111000"
        )
    port map (
            in0 => \N__5912\,
            in1 => \N__6628\,
            in2 => \N__5984\,
            in3 => \N__6738\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0\,
            ltout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_2_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__5970\,
            in1 => \N__6635\,
            in2 => \N__5957\,
            in3 => \N__5952\,
            lcout => \U712_CHIP_RAM.SDRAM_CMDZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9719\,
            ce => \N__5936\,
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_2_0_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111001010"
        )
    port map (
            in0 => \N__6619\,
            in1 => \N__5908\,
            in2 => \N__6222\,
            in3 => \N__6734\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.N_316_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_1_0_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110100"
        )
    port map (
            in0 => \N__6735\,
            in1 => \N__6211\,
            in2 => \N__6644\,
            in3 => \N__6408\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_2_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110110101000"
        )
    port map (
            in0 => \N__6214\,
            in1 => \N__6496\,
            in2 => \N__6416\,
            in3 => \N__6621\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_0_101_i_a2_0_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_3_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110100101000"
        )
    port map (
            in0 => \N__6213\,
            in1 => \N__6495\,
            in2 => \N__6415\,
            in3 => \N__6620\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_138_i_a2_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNO_0_0_LC_10_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__6494\,
            in2 => \_gnd_net_\,
            in3 => \N__6407\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_cnst_0_2_29_i_a2_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_CYCLE_START_RNIBRI34_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__6299\,
            in1 => \N__6223\,
            in2 => \_gnd_net_\,
            in3 => \N__6097\,
            lcout => \U712_CHIP_RAM.N_109_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_TACK_RNO_1_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6780\,
            in1 => \N__6835\,
            in2 => \_gnd_net_\,
            in3 => \N__7206\,
            lcout => \U712_REG_SM.un15_0_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNIELLV_7_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__7205\,
            in1 => \N__8319\,
            in2 => \_gnd_net_\,
            in3 => \N__8251\,
            lcout => \U712_REG_SM.LATCH_REG_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__8083\,
            in1 => \N__10879\,
            in2 => \_gnd_net_\,
            in3 => \N__6904\,
            lcout => \REG_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.REG_TACK_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000111100000"
        )
    port map (
            in0 => \N__6905\,
            in1 => \N__6896\,
            in2 => \N__6890\,
            in3 => \N__6865\,
            lcout => \REG_TACK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.C1_SYNC_1_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7481\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.STATE_COUNTER_7_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011101010"
        )
    port map (
            in0 => \N__6836\,
            in1 => \N__8326\,
            in2 => \N__7213\,
            in3 => \N__8259\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.C3_SYNC_1_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7109\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.REGENn_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__6811\,
            in1 => \N__7957\,
            in2 => \_gnd_net_\,
            in3 => \N__8084\,
            lcout => \REGENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.STATE_COUNTER_4_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6784\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.STATE_COUNTER_3_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8378\,
            in1 => \N__8327\,
            in2 => \N__8261\,
            in3 => \N__6760\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLEC_net\,
            ce => 'H',
            sr => \N__10976\
        );

    \U712_REG_SM.STATE_COUNTER_2_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111010000"
        )
    port map (
            in0 => \N__6764\,
            in1 => \N__7178\,
            in2 => \N__8392\,
            in3 => \N__7961\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.STATE_COUNTER_2C_net\,
            ce => 'H',
            sr => \N__10974\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_5_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111010101"
        )
    port map (
            in0 => \N__8634\,
            in1 => \N__7097\,
            in2 => \N__10692\,
            in3 => \N__9569\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_1_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10686\,
            in1 => \N__7103\,
            in2 => \N__9137\,
            in3 => \N__8120\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_5_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8633\,
            in1 => \N__7096\,
            in2 => \N__10693\,
            in3 => \N__9568\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_7_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10639\,
            in1 => \N__7073\,
            in2 => \N__9136\,
            in3 => \N__7061\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI4VDC_0_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9172\,
            in2 => \_gnd_net_\,
            in3 => \N__8915\,
            lcout => \U712_CHIP_RAM.CMA_5_sn_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9617\,
            in1 => \N__9554\,
            in2 => \_gnd_net_\,
            in3 => \N__9968\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_3C_net\,
            ce => \N__9773\,
            sr => \N__10994\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9969\,
            in1 => \N__9485\,
            in2 => \_gnd_net_\,
            in3 => \N__9406\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_7C_net\,
            ce => \N__9770\,
            sr => \N__10989\
        );

    \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__7039\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7008\,
            lcout => \U712_BYTE_ENABLE.un1_CUMBEn_i_0_a3_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_0_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__7768\,
            in1 => \N__7783\,
            in2 => \N__7754\,
            in3 => \N__7798\,
            lcout => \U712_CHIP_RAM.REFRESH5lt7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_49_i_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110111011101"
        )
    port map (
            in0 => \N__6944\,
            in1 => \N__10837\,
            in2 => \N__7250\,
            in3 => \N__10647\,
            lcout => \N_49_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.LMBE_i_o4_0_o3_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000111011"
        )
    port map (
            in0 => \N__10347\,
            in1 => \N__10251\,
            in2 => \N__10181\,
            in3 => \N__10407\,
            lcout => \U712_BYTE_ENABLE.N_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BUFFERS.DRDDIR_0_m2_i_m2_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001111111"
        )
    port map (
            in0 => \N__10775\,
            in1 => \N__10864\,
            in2 => \N__7926\,
            in3 => \N__7426\,
            lcout => \N_315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIGHT91_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__8250\,
            in2 => \N__8282\,
            in3 => \N__7204\,
            lcout => \U712_REG_SM.N_278\,
            ltout => \U712_REG_SM.N_278_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C1_SYNC_RNI5ITS1_1_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111010"
        )
    port map (
            in0 => \N__8398\,
            in1 => \_gnd_net_\,
            in2 => \N__7217\,
            in3 => \N__8318\,
            lcout => \U712_REG_SM.C1_SYNC_RNI5ITS1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_1_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__7174\,
            in1 => \N__7162\,
            in2 => \N__8399\,
            in3 => \N__8421\,
            lcout => \U712_REG_SM.UDSn_7_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.STATE_COUNTER_RNI5J3V_7_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__8479\,
            in1 => \N__7919\,
            in2 => \_gnd_net_\,
            in3 => \N__7203\,
            lcout => \U712_REG_SM.N_309\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_RNI6FIN_1_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__8249\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8317\,
            lcout => \U712_REG_SM.N_272\,
            ltout => \U712_REG_SM.N_272_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_1_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__7163\,
            in1 => \N__8394\,
            in2 => \N__7154\,
            in3 => \N__7335\,
            lcout => \U712_REG_SM.LDSn_7_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.C3_SYNC_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7132\,
            lcout => \U712_REG_SM.C3_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10975\
        );

    \U712_REG_SM.C1_SYNC_0_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7517\,
            lcout => \U712_REG_SM.C1_SYNCZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10975\
        );

    \U712_REG_SM.LDSn_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__7310\,
            in1 => \N__7336\,
            in2 => \N__7475\,
            in3 => \N__7634\,
            lcout => \LDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10975\
        );

    \U712_REG_SM.ASn_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__7463\,
            in1 => \N__7441\,
            in2 => \N__8336\,
            in3 => \N__8085\,
            lcout => \ASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.C3_SYNC_0C_net\,
            ce => 'H',
            sr => \N__10975\
        );

    \U712_BUFFERS.DMA_LATCH_EN_i_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000111"
        )
    port map (
            in0 => \N__10857\,
            in1 => \N__10763\,
            in2 => \N__7430\,
            in3 => \N__7873\,
            lcout => \N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_2_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7334\,
            in2 => \_gnd_net_\,
            in3 => \N__8375\,
            lcout => OPEN,
            ltout => \U712_REG_SM.N_467_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.LDSn_RNO_0_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000000"
        )
    port map (
            in0 => \N__10130\,
            in1 => \N__10259\,
            in2 => \N__7313\,
            in3 => \N__8491\,
            lcout => \U712_REG_SM.N_371\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_1_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7616\,
            in1 => \N__7622\,
            in2 => \_gnd_net_\,
            in3 => \N__7304\,
            lcout => \CMA_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9714\,
            ce => \N__9647\,
            sr => \N__10999\
        );

    \U712_CHIP_RAM.CMA_esr_5_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__7289\,
            in1 => \N__7283\,
            in2 => \_gnd_net_\,
            in3 => \N__7256\,
            lcout => \CMA_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9714\,
            ce => \N__9647\,
            sr => \N__10999\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_5_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__8750\,
            in1 => \N__9118\,
            in2 => \_gnd_net_\,
            in3 => \N__7586\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_1_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001011110000"
        )
    port map (
            in0 => \N__8584\,
            in1 => \N__10641\,
            in2 => \N__8773\,
            in3 => \N__9117\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_2_1_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111011111111"
        )
    port map (
            in0 => \N__8585\,
            in1 => \N__10640\,
            in2 => \N__8774\,
            in3 => \N__9116\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_2_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__7610\,
            in1 => \N__10655\,
            in2 => \N__9122\,
            in3 => \N__7535\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_0_3_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__8919\,
            in1 => \N__9173\,
            in2 => \N__8972\,
            in3 => \N__9090\,
            lcout => \U712_CHIP_RAM.REFRESH_RST\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_3_5_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__7601\,
            in1 => \N__10654\,
            in2 => \N__8102\,
            in3 => \_gnd_net_\,
            lcout => \U712_CHIP_RAM.N_329\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_1_0_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__7580\,
            in1 => \N__7562\,
            in2 => \_gnd_net_\,
            in3 => \N__9076\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_1Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.REFRESH_RNO_1_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7718\,
            in2 => \_gnd_net_\,
            in3 => \N__7736\,
            lcout => \U712_CHIP_RAM.REFRESH5lto7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9537\,
            in1 => \N__10076\,
            in2 => \_gnd_net_\,
            in3 => \N__9961\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_2C_net\,
            ce => \N__9771\,
            sr => \N__10981\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7526\,
            in2 => \_gnd_net_\,
            in3 => \N__7520\,
            lcout => \U712_CHIP_RAM.REFRESH5lto0\,
            ltout => OPEN,
            carryin => \bfn_12_10_0_\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7799\,
            in2 => \_gnd_net_\,
            in3 => \N__7787\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_0\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_2_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7784\,
            in2 => \_gnd_net_\,
            in3 => \N__7772\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_2\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_1\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7769\,
            in2 => \_gnd_net_\,
            in3 => \N__7757\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_3\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_2\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_4_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7753\,
            in2 => \_gnd_net_\,
            in3 => \N__7739\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_4\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_3\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_5_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7735\,
            in2 => \_gnd_net_\,
            in3 => \N__7721\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_5\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_4\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_6_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7717\,
            in2 => \_gnd_net_\,
            in3 => \N__7703\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_6\,
            ltout => OPEN,
            carryin => \U712_CHIP_RAM.REFRESH_COUNTER_cry_5\,
            carryout => \U712_CHIP_RAM.REFRESH_COUNTER_cry_6\,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_CHIP_RAM.REFRESH_COUNTER_7_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7693\,
            in2 => \_gnd_net_\,
            in3 => \N__7700\,
            lcout => \U712_CHIP_RAM.REFRESH_COUNTERZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__7674\,
            ce => 'H',
            sr => \N__7652\
        );

    \U712_REG_SM.UDSn_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__7640\,
            in1 => \N__8447\,
            in2 => \N__8428\,
            in3 => \N__7633\,
            lcout => \UDSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10973\
        );

    \U712_REG_SM.STATE_COUNTER_0_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__8086\,
            in1 => \N__8216\,
            in2 => \_gnd_net_\,
            in3 => \N__8490\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.UDSnC_net\,
            ce => 'H',
            sr => \N__10973\
        );

    \U712_REG_SM.REG_CYCLE_START_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011011100000101"
        )
    port map (
            in0 => \N__8044\,
            in1 => \N__7970\,
            in2 => \N__8012\,
            in3 => \N__8281\,
            lcout => \U712_REG_SM.REG_CYCLE_STARTZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \N__10972\
        );

    \U712_REG_SM.CYCLE_RUN_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011100"
        )
    port map (
            in0 => \N__8214\,
            in1 => \N__7969\,
            in2 => \N__8492\,
            in3 => \N__7950\,
            lcout => \U712_REG_SM.CYCLE_RUNZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \N__10972\
        );

    \U712_REG_SM.STATE_COUNTER_1_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8213\,
            in2 => \_gnd_net_\,
            in3 => \N__8488\,
            lcout => \U712_REG_SM.STATE_COUNTERZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \N__10972\
        );

    \U712_REG_SM.REG_WRITE_CYCLE_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111000001110100"
        )
    port map (
            in0 => \N__7927\,
            in1 => \N__8489\,
            in2 => \N__7879\,
            in3 => \N__8215\,
            lcout => \REG_WRITE_CYCLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_REG_SM.REG_CYCLE_STARTC_net\,
            ce => 'H',
            sr => \N__10972\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNIA0SO_3_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__9183\,
            in1 => \N__9123\,
            in2 => \N__8980\,
            in3 => \N__8928\,
            lcout => OPEN,
            ltout => \U712_CHIP_RAM.un1_CMA28_0_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI0AO81_3_LC_13_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__7844\,
            in3 => \N__11030\,
            lcout => \U712_CHIP_RAM.un1_CMA28_0_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8775\,
            in1 => \N__8594\,
            in2 => \N__8726\,
            in3 => \N__8144\,
            lcout => \CMA_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9716\,
            ce => \N__9655\,
            sr => \N__11002\
        );

    \U712_CHIP_RAM.CMA_esr_2_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8776\,
            in1 => \N__9812\,
            in2 => \N__8727\,
            in3 => \N__7823\,
            lcout => \CMA_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9716\,
            ce => \N__9655\,
            sr => \N__11002\
        );

    \U712_CHIP_RAM.CMA_esr_7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8777\,
            in1 => \N__8718\,
            in2 => \N__9437\,
            in3 => \N__8180\,
            lcout => \CMA_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9716\,
            ce => \N__9655\,
            sr => \N__11002\
        );

    \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9_1_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9124\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \U712_CHIP_RAM.SDRAM_CMD_RNI8NM9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_0_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10671\,
            in1 => \N__8150\,
            in2 => \N__9138\,
            in3 => \N__8573\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_6_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101000"
        )
    port map (
            in0 => \N__8138\,
            in1 => \N__10673\,
            in2 => \N__9140\,
            in3 => \N__8093\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CMA_esr_RNO_0_4_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111001000"
        )
    port map (
            in0 => \N__10672\,
            in1 => \N__8129\,
            in2 => \N__9139\,
            in3 => \N__8108\,
            lcout => \U712_CHIP_RAM.CMA_esr_RNO_0Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1_LC_13_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10075\,
            in1 => \N__10023\,
            in2 => \_gnd_net_\,
            in3 => \N__9948\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9775\,
            sr => \N__10990\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_4_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9358\,
            in1 => \N__9611\,
            in2 => \_gnd_net_\,
            in3 => \N__9949\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9775\,
            sr => \N__10990\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_5_LC_13_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9950\,
            in1 => \N__9359\,
            in2 => \_gnd_net_\,
            in3 => \N__9325\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9775\,
            sr => \N__10990\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_6_LC_13_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9326\,
            in1 => \N__9484\,
            in2 => \_gnd_net_\,
            in3 => \N__9951\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_1C_net\,
            ce => \N__9775\,
            sr => \N__10990\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_0_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9959\,
            in1 => \N__8528\,
            in2 => \_gnd_net_\,
            in3 => \N__8556\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9798\,
            ce => \N__9774\,
            sr => \N__10983\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_1_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9960\,
            in1 => \N__8557\,
            in2 => \_gnd_net_\,
            in3 => \N__10025\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9798\,
            ce => \N__9774\,
            sr => \N__10983\
        );

    \U712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__8564\,
            in1 => \N__10019\,
            in2 => \_gnd_net_\,
            in3 => \N__9933\,
            lcout => \U712_CHIP_RAM.DMA_COL_ADDRESSZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9772\,
            sr => \N__10982\
        );

    \U712_CHIP_RAM.DMA_A1_nesr_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__8563\,
            in1 => \N__8521\,
            in2 => \_gnd_net_\,
            in3 => \N__9932\,
            lcout => \U712_CHIP_RAM.DMA_AZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVU712_CHIP_RAM.DMA_COL_ADDRESS_nesr_0C_net\,
            ce => \N__9772\,
            sr => \N__10982\
        );

    \U712_REG_SM.UDSn_RNO_0_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__10281\,
            in1 => \N__8342\,
            in2 => \N__10187\,
            in3 => \N__8484\,
            lcout => \U712_REG_SM.N_369\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.UDSn_RNO_2_LC_13_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8420\,
            in2 => \_gnd_net_\,
            in3 => \N__8393\,
            lcout => \U712_REG_SM.N_465\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_REG_SM.REG_CYCLE_START_RNIPBK41_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__8331\,
            in1 => \N__8280\,
            in2 => \_gnd_net_\,
            in3 => \N__8260\,
            lcout => \U712_REG_SM.N_288\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.CASn_LC_14_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9135\,
            lcout => \CASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9713\,
            ce => 'H',
            sr => \N__11014\
        );

    \U712_CHIP_RAM.WEn_LC_14_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8935\,
            lcout => \WEn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9713\,
            ce => 'H',
            sr => \N__11014\
        );

    \U712_CHIP_RAM.RASn_LC_14_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9191\,
            lcout => \RASn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9713\,
            ce => 'H',
            sr => \N__11014\
        );

    \U712_CHIP_RAM.CRCSn_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8979\,
            lcout => \CRCSn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9715\,
            ce => 'H',
            sr => \N__11013\
        );

    \U712_CHIP_RAM.CMA_esr_10_LC_14_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__9190\,
            in1 => \N__9134\,
            in2 => \N__8981\,
            in3 => \N__8936\,
            lcout => \CMA_c_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9717\,
            ce => \N__9654\,
            sr => \N__11012\
        );

    \U712_CHIP_RAM.CMA_esr_8_LC_14_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__8645\,
            in1 => \N__8873\,
            in2 => \N__10697\,
            in3 => \N__9494\,
            lcout => \CMA_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9717\,
            ce => \N__9654\,
            sr => \N__11012\
        );

    \U712_CHIP_RAM.CMA_esr_3_LC_14_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8778\,
            in1 => \N__9503\,
            in2 => \N__8728\,
            in3 => \N__8831\,
            lcout => \CMA_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9718\,
            ce => \N__9659\,
            sr => \N__11007\
        );

    \U712_CHIP_RAM.CMA_esr_6_LC_14_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__8780\,
            in1 => \N__8725\,
            in2 => \N__9281\,
            in3 => \N__8807\,
            lcout => \CMA_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9718\,
            ce => \N__9659\,
            sr => \N__11007\
        );

    \U712_CHIP_RAM.CMA_esr_4_LC_14_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__8779\,
            in1 => \N__9623\,
            in2 => \N__8729\,
            in3 => \N__8693\,
            lcout => \CMA_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9718\,
            ce => \N__9659\,
            sr => \N__11007\
        );

    \U712_CHIP_RAM.CMA_esr_9_LC_14_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000110010000000"
        )
    port map (
            in0 => \N__8666\,
            in1 => \N__8641\,
            in2 => \N__10691\,
            in3 => \N__9368\,
            lcout => \CMA_c_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9718\,
            ce => \N__9659\,
            sr => \N__11007\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_4_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__9553\,
            in1 => \N__9612\,
            in2 => \_gnd_net_\,
            in3 => \N__9924\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9800\,
            ce => \N__9778\,
            sr => \N__11003\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_5_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__9357\,
            in1 => \N__9613\,
            in2 => \_gnd_net_\,
            in3 => \N__9925\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9800\,
            ce => \N__9778\,
            sr => \N__11003\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_3_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__10067\,
            in1 => \N__9546\,
            in2 => \_gnd_net_\,
            in3 => \N__9908\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => \N__9777\,
            sr => \N__10995\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_8_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9910\,
            in1 => \N__9477\,
            in2 => \_gnd_net_\,
            in3 => \N__9398\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => \N__9777\,
            sr => \N__10995\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_7_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9909\,
            in1 => \N__9324\,
            in2 => \_gnd_net_\,
            in3 => \N__9476\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => \N__9777\,
            sr => \N__10995\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_9_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__9911\,
            in1 => \N__9425\,
            in2 => \_gnd_net_\,
            in3 => \N__9399\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9799\,
            ce => \N__9777\,
            sr => \N__10995\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_6_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__9907\,
            in1 => \N__9351\,
            in2 => \_gnd_net_\,
            in3 => \N__9323\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9797\,
            ce => \N__9776\,
            sr => \N__10991\
        );

    \U712_BYTE_ENABLE.N_50_i_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000111110011"
        )
    port map (
            in0 => \N__10475\,
            in1 => \N__10516\,
            in2 => \N__10782\,
            in3 => \N__10678\,
            lcout => \N_50_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UUBE_i_o4_0_o3_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001111010111"
        )
    port map (
            in0 => \N__10186\,
            in1 => \N__10258\,
            in2 => \N__10423\,
            in3 => \N__10349\,
            lcout => OPEN,
            ltout => \U712_BYTE_ENABLE.N_91_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_51_i_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__10679\,
            in1 => \N__10517\,
            in2 => \N__10499\,
            in3 => \N__10836\,
            lcout => \N_51_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.UMBE_i_o4_0_o3_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101011111000111"
        )
    port map (
            in0 => \N__10348\,
            in1 => \N__10416\,
            in2 => \N__10272\,
            in3 => \N__10185\,
            lcout => \U712_BYTE_ENABLE.N_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_90_i_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101001100"
        )
    port map (
            in0 => \N__10336\,
            in1 => \N__10276\,
            in2 => \N__10179\,
            in3 => \N__10404\,
            lcout => \N_90_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_92_i_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101000010010"
        )
    port map (
            in0 => \N__10406\,
            in1 => \N__10338\,
            in2 => \N__10283\,
            in3 => \N__10167\,
            lcout => \N_92_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_91_i_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001011001000"
        )
    port map (
            in0 => \N__10337\,
            in1 => \N__10277\,
            in2 => \N__10180\,
            in3 => \N__10405\,
            lcout => \N_91_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_BYTE_ENABLE.N_89_i_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100001011000"
        )
    port map (
            in0 => \N__10403\,
            in1 => \N__10335\,
            in2 => \N__10282\,
            in3 => \N__10160\,
            lcout => \N_89_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \U712_CHIP_RAM.DMA_ROW_ADDRESS_esr_2_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__10068\,
            in1 => \N__10024\,
            in2 => \_gnd_net_\,
            in3 => \N__9955\,
            lcout => \U712_CHIP_RAM.DMA_ROW_ADDRESSZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__9796\,
            ce => \N__9779\,
            sr => \N__11008\
        );

    \U712_BUFFERS.un1_DRDENn_LC_24_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__10895\,
            in1 => \N__10832\,
            in2 => \_gnd_net_\,
            in3 => \N__10740\,
            lcout => \DRDENn_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
